* NGSPICE file created from team_05_Wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_16 abstract view
.subckt sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

.subckt team_05_Wrapper ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14]
+ ADR_O[15] ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22]
+ ADR_O[23] ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30]
+ ADR_O[31] ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0]
+ DAT_I[10] DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17]
+ DAT_I[18] DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25]
+ DAT_I[26] DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4]
+ DAT_I[5] DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12]
+ DAT_O[13] DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20]
+ DAT_O[21] DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28]
+ DAT_O[29] DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7]
+ DAT_O[8] DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[34] gpio_in[35] gpio_in[36]
+ gpio_in[37] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9]
+ gpio_oeb[0] gpio_oeb[10] gpio_oeb[11] gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15]
+ gpio_oeb[16] gpio_oeb[17] gpio_oeb[18] gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21]
+ gpio_oeb[22] gpio_oeb[23] gpio_oeb[24] gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28]
+ gpio_oeb[29] gpio_oeb[2] gpio_oeb[30] gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[34]
+ gpio_oeb[35] gpio_oeb[36] gpio_oeb[37] gpio_oeb[3] gpio_oeb[4] gpio_oeb[5] gpio_oeb[6]
+ gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12]
+ gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19]
+ gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25]
+ gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31]
+ gpio_out[32] gpio_out[33] gpio_out[34] gpio_out[35] gpio_out[36] gpio_out[37] gpio_out[3]
+ gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] irq[0] irq[1]
+ irq[2] la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13]
+ la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19]
+ la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24]
+ la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2]
+ la_data_in[30] la_data_in[31] la_data_in[3] la_data_in[4] la_data_in[5] la_data_in[6]
+ la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10] la_data_out[11]
+ la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16]
+ la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21]
+ la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26]
+ la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31]
+ la_data_out[3] la_data_out[4] la_data_out[5] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[3] la_oenb[4]
+ la_oenb[5] la_oenb[6] la_oenb[7] la_oenb[8] la_oenb[9] vccd1 vssd1 wb_clk_i wb_rst_i
+ wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XANTENNA__09523__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09671_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[1\]
+ net876 net874 net860 vssd1 vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__and4_1
XANTENNA__08731__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08622_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[24\]
+ net717 _04691_ _04696_ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__o22ai_1
XANTENNA__13607__A1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11618__B1 _07472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08553_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[26\]
+ net824 net784 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[26\]
+ _04619_ vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08484_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[27\]
+ net692 net599 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18363__1348 vssd1 vssd1 vccd1 vccd1 _18363__1348/HI net1348 sky130_fd_sc_hd__conb_1
XFILLER_0_58_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1071_A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout427_A _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1169_A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08798__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09105_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[12\]
+ net660 _05161_ net719 vssd1 vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__a211o_1
XFILLER_0_73_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout215_X net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09036_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[14\]
+ net775 net765 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[14\]
+ _05095_ vssd1 vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__a221o_1
XFILLER_0_130_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout796_A net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13496__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold340 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[37\] vssd1 vssd1
+ vccd1 vccd1 net1754 sky130_fd_sc_hd__dlygate4sd3_1
Xhold351 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[67\] vssd1 vssd1
+ vccd1 vccd1 net1765 sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[100\] vssd1 vssd1
+ vccd1 vccd1 net1776 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold373 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[51\] vssd1 vssd1
+ vccd1 vccd1 net1787 sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[27\] vssd1 vssd1
+ vccd1 vccd1 net1798 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09762__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold395 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[4\] vssd1 vssd1
+ vccd1 vccd1 net1809 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout963_A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09706__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout820 net821 vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__clkbuf_4
Xfanout831 net832 vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__buf_4
XFILLER_0_102_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09938_ _05935_ _05936_ vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__or2_1
Xfanout842 net844 vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__clkbuf_8
Xfanout853 _04367_ vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__clkbuf_8
Xfanout864 net866 vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__buf_2
Xfanout875 _04283_ vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout886 _04281_ vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__buf_2
X_09869_ _05897_ vssd1 vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__inv_2
Xfanout897 net898 vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__buf_4
XANTENNA_fanout751_X net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1040 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2454 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11321__A2 _07097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17642__D team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1051 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2465 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08722__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout849_X net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1062 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2476 sky130_fd_sc_hd__dlygate4sd3_1
X_11900_ _07676_ _07711_ _07677_ vssd1 vssd1 vccd1 vccd1 _07712_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09722__B net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12880_ net283 net2805 net479 vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__mux2_1
Xhold1073 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1084 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 net2498 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1095 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 net2509 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _07590_ _07629_ _07640_ vssd1 vssd1 vccd1 vccd1 _07643_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_159_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_159_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ net1084 vssd1 vssd1 vccd1 vccd1 _00180_ sky130_fd_sc_hd__inv_2
X_11762_ _07531_ _07558_ vssd1 vssd1 vccd1 vccd1 _07574_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13501_ net2605 net235 net405 vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10713_ _05597_ net553 net334 _06252_ _06713_ vssd1 vssd1 vccd1 vccd1 _06714_ sky130_fd_sc_hd__o221a_1
XANTENNA__12575__S net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14481_ net1188 vssd1 vssd1 vccd1 vccd1 _00111_ sky130_fd_sc_hd__inv_2
X_11693_ team_05_WB.EN_VAL_REG net72 _07505_ vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16220_ net1090 vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__inv_2
XANTENNA__12034__B1 _07352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13432_ net2922 net223 net414 vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__mux2_1
X_10644_ _05577_ _06017_ _06049_ _06644_ vssd1 vssd1 vccd1 vccd1 _06649_ sky130_fd_sc_hd__o31a_1
XFILLER_0_125_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16151_ net1153 vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__inv_2
X_10575_ _05826_ net511 _06263_ _06510_ _06577_ vssd1 vssd1 vccd1 vccd1 _06584_ sky130_fd_sc_hd__o221a_1
X_13363_ net2014 net194 net421 vssd1 vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__mux2_1
XANTENNA__08253__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15102_ net1066 vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__inv_2
X_12314_ _03542_ net251 _03602_ vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__a21o_1
X_16082_ net1174 vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__inv_2
XANTENNA__08641__X team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[24\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13294_ net307 net2760 net432 vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__mux2_1
XANTENNA__15187__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15033_ net1052 vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12245_ _03510_ _03539_ _03538_ _03537_ vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_122_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12176_ _07933_ _07937_ _07938_ _07941_ vssd1 vssd1 vccd1 vccd1 _07988_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_20_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09616__C net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11127_ _07058_ _07052_ vssd1 vssd1 vccd1 vccd1 _07093_ sky130_fd_sc_hd__and2b_2
X_16984_ clknet_leaf_32_wb_clk_i _02614_ _00680_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11058_ _07023_ _07024_ vssd1 vssd1 vccd1 vccd1 _07025_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15935_ net1300 vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__inv_2
XANTENNA__09505__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_60_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11312__A2 _07117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08713__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10009_ _04989_ net365 vssd1 vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__or2_1
X_15866_ net1290 vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__inv_2
XANTENNA__09632__B net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10520__B1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17605_ clknet_leaf_81_wb_clk_i _02976_ _01301_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_14817_ net1236 vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__inv_2
X_15797_ net1297 vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__inv_2
X_17536_ clknet_leaf_81_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[7\]
+ _01232_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14748_ net1063 vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_48_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_80_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12485__S net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17467_ clknet_leaf_38_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[2\]
+ _01163_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08492__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14679_ net1099 vssd1 vssd1 vccd1 vccd1 _00309_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16418_ clknet_leaf_6_wb_clk_i _02048_ _00114_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17398_ clknet_leaf_59_wb_clk_i net1426 _01094_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_172_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16349_ clknet_leaf_109_wb_clk_i _01979_ _00045_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08244__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14317__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[19\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18019_ clknet_leaf_96_wb_clk_i _03358_ _01715_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10339__A0 _06060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09723_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[0\]
+ net944 net1014 net934 vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__and4_1
XANTENNA_clkbuf_leaf_87_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_59_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09654_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[1\]
+ net829 _05676_ _05681_ _05685_ vssd1 vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_87_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08605_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[24\]
+ net634 net618 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_26_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_943 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09585_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[2\]
+ net948 net933 net930 vssd1 vssd1 vccd1 vccd1 _05621_ sky130_fd_sc_hd__and4_1
XFILLER_0_139_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1286_A net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08536_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[26\]
+ net718 _04609_ _04612_ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_166_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12395__S _03660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout332_X net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout711_A _04288_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08467_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[28\]
+ net828 _04545_ net856 vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__a211o_1
XANTENNA__08483__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09417__D1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08398_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[29\]
+ net700 net624 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__a22o_1
XANTENNA__12567__A1 _07797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13764__B1 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10578__B1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1241_X net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10360_ _06063_ _06379_ _06375_ _06371_ vssd1 vssd1 vccd1 vccd1 _06380_ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17637__D team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout799_X net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09019_ _04355_ _05079_ vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__nand2_1
X_10291_ _06100_ _06313_ vssd1 vssd1 vccd1 vccd1 _06314_ sky130_fd_sc_hd__or2_1
XANTENNA__09717__B net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12030_ _07369_ _07841_ vssd1 vssd1 vccd1 vccd1 _07842_ sky130_fd_sc_hd__or2_1
XANTENNA__09196__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold170 net90 vssd1 vssd1 vccd1 vccd1 net1584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[6\]
+ vssd1 vssd1 vccd1 vccd1 net1595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 net129 vssd1 vssd1 vccd1 vccd1 net1606 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08943__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08340__C _04418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout650 net651 vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_109_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout661 net662 vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11982__B _07791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout672 net675 vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__buf_6
X_13981_ _03828_ _03831_ _03851_ vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__or3b_1
Xfanout683 net686 vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__clkbuf_8
Xfanout694 _04297_ vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__buf_4
X_15720_ net1142 vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__inv_2
X_12932_ net191 net2471 net469 vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_126_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10598__B _06605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15651_ net1250 vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__inv_2
X_12863_ net193 net2784 net477 vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__mux2_1
X_14602_ net1110 vssd1 vssd1 vccd1 vccd1 _00232_ sky130_fd_sc_hd__inv_2
X_18370_ net1355 vssd1 vssd1 vccd1 vccd1 la_data_out[18] sky130_fd_sc_hd__buf_2
X_11814_ _07605_ _07609_ _07598_ _07599_ vssd1 vssd1 vccd1 vccd1 _07626_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_157_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15582_ net1251 vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12794_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[10\] _04255_
+ vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_164_Left_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09120__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17321_ clknet_leaf_21_wb_clk_i _02951_ _01017_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_174_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ net1191 vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_174_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13702__B _06729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11745_ _07546_ _07556_ _07540_ vssd1 vssd1 vccd1 vccd1 _07557_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17252_ clknet_leaf_193_wb_clk_i _02882_ _00948_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14464_ net1200 vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__inv_2
X_11676_ _07488_ _07490_ team_05_WB.instance_to_wrap.wishbone.curr_state\[0\] vssd1
+ vssd1 vccd1 vccd1 _07491_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_12_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16203_ net1072 vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13415_ net2834 net291 net416 vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__mux2_1
X_10627_ _06338_ _06510_ _06630_ _06631_ _06632_ vssd1 vssd1 vccd1 vccd1 _06633_ sky130_fd_sc_hd__o2111a_1
X_17183_ clknet_leaf_152_wb_clk_i _02813_ _00879_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14395_ net1506 vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10569__B1 _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16134_ net1306 vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13346_ net277 net2856 net427 vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__mux2_1
X_10558_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[12\] _06091_ vssd1
+ vssd1 vccd1 vccd1 _06568_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16065_ net1173 vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13277_ net259 net2869 net432 vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__mux2_1
X_10489_ _06500_ _06501_ net892 vssd1 vssd1 vccd1 vccd1 _06502_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09187__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_173_Left_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15016_ net1224 vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__inv_2
X_12228_ _03521_ _03522_ vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__or2_1
XANTENNA__09726__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_121_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_166_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08934__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12159_ _07919_ _07969_ vssd1 vssd1 vccd1 vccd1 _07971_ sky130_fd_sc_hd__xnor2_1
X_18362__1347 vssd1 vssd1 vccd1 vccd1 _18362__1347/HI net1347 sky130_fd_sc_hd__conb_1
XFILLER_0_75_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16967_ clknet_leaf_201_wb_clk_i _02597_ _00663_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15918_ net1267 vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__inv_2
X_16898_ clknet_leaf_3_wb_clk_i _02528_ _00594_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15849_ net1273 vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09370_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[7\]
+ net816 net788 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[7\]
+ _05402_ vssd1 vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_82_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09111__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10257__C1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08321_ net942 net931 net928 vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17519_ clknet_leaf_73_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[22\]
+ _01215_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08465__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13104__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08252_ _04328_ _04330_ _04332_ _04334_ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__or4_1
XFILLER_0_7_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12549__A1 _07789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08183_ _04231_ _04237_ vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__nor2_1
XANTENNA__12943__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_160_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10029__A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08281__X _04363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1034_A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09178__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_15__f_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout494_A _03699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_89_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout661_A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout282_X net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09706_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[0\]
+ net945 net936 net934 vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__and4_1
XFILLER_0_156_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08169__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09637_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[1\]
+ net1015 net940 net924 vssd1 vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__and4_1
XFILLER_0_97_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09568_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[2\]
+ net946 net939 _04418_ vssd1 vssd1 vccd1 vccd1 _05604_ sky130_fd_sc_hd__and4_1
XFILLER_0_167_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09102__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08519_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[26\]
+ net702 net609 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__a22o_1
X_09499_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[4\]
+ net680 net630 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[4\]
+ _05537_ vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout714_X net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08456__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13014__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11530_ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[28\] _07440_ _07345_
+ vssd1 vssd1 vccd1 vccd1 _07441_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08335__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_137_Right_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11461_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[7\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[7\]
+ net1034 vssd1 vssd1 vccd1 vccd1 _07372_ sky130_fd_sc_hd__mux2_1
XANTENNA__12853__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08208__A2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13200_ _06317_ net2729 net352 vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__mux2_1
X_10412_ _06034_ _06044_ vssd1 vssd1 vccd1 vccd1 _06429_ sky130_fd_sc_hd__nand2_1
X_11392_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[5\] _07322_
+ vssd1 vssd1 vccd1 vccd1 _07323_ sky130_fd_sc_hd__and2_1
X_14180_ team_05_WB.instance_to_wrap.CPU_DAT_O\[29\] net504 net908 vssd1 vssd1 vccd1
+ vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[29\] sky130_fd_sc_hd__and3_1
XFILLER_0_33_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13131_ net220 net2258 net446 vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__mux2_1
X_10343_ _06099_ _06363_ vssd1 vssd1 vccd1 vccd1 _06364_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09169__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input55_A wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10274_ net555 _06296_ vssd1 vssd1 vccd1 vccd1 _06297_ sky130_fd_sc_hd__nor2_1
X_13062_ net199 net2719 net454 vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13684__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08916__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12013_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[30\] team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[15\]
+ net995 net548 vssd1 vssd1 vccd1 vccd1 _07825_ sky130_fd_sc_hd__a31o_1
X_17870_ clknet_leaf_76_wb_clk_i _03213_ _01566_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[52\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16821_ clknet_leaf_24_wb_clk_i _02451_ _00517_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout480 net483 vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_6_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout491 _03700_ vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__clkbuf_4
X_16752_ clknet_leaf_151_wb_clk_i _02382_ _00448_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13964_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[3\] _03805_ _03836_
+ _07451_ vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__o211a_1
XANTENNA__09613__D net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15703_ net1166 vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__inv_2
XANTENNA__09341__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12915_ net292 net2436 net472 vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__mux2_1
X_16683_ clknet_leaf_188_wb_clk_i _02313_ _00379_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13895_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[19\]
+ net558 net574 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[19\]
+ net985 vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__a221o_1
XANTENNA__08695__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13713__A net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15634_ net1282 vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12846_ net275 net2758 net482 vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08807__A net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18353_ net1338 vssd1 vssd1 vccd1 vccd1 la_data_out[1] sky130_fd_sc_hd__buf_2
X_15565_ net1246 vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12777_ net271 net2705 net488 vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__mux2_1
XANTENNA__08447__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17304_ clknet_leaf_28_wb_clk_i _02934_ _01000_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14516_ net1073 vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__inv_2
X_18284_ net107 vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__clkbuf_1
X_11728_ _07534_ _07539_ vssd1 vssd1 vccd1 vccd1 _07540_ sky130_fd_sc_hd__nor2_1
X_15496_ net1159 vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17235_ clknet_leaf_167_wb_clk_i _02865_ _00931_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14447_ net1233 vssd1 vssd1 vccd1 vccd1 _00077_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11659_ net3 net992 _07483_ net1642 vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__a22o_1
XANTENNA__12763__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11203__A1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17166_ clknet_leaf_170_wb_clk_i _02796_ _00862_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14378_ net1540 vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold906 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net2320 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11379__S net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16117_ net1134 vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__inv_2
Xhold917 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2331 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13329_ net199 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[31\]
+ net426 vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__mux2_1
Xhold928 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold939 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17097_ clknet_leaf_21_wb_clk_i _02727_ _00793_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16048_ net1251 vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08907__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13594__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12351__X _03646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08870_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[17\]
+ net707 net679 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_32_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17999_ clknet_leaf_63_wb_clk_i _03338_ _01695_ vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_84_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09332__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12938__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08686__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09422_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[5\]
+ net714 net641 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05465_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13967__B1 _07451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09353_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[27\] _04246_
+ _04350_ _05399_ vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__o31a_1
XANTENNA__08438__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08304_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[31\]
+ net834 net830 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[31\]
+ _04385_ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__a221o_1
XFILLER_0_142_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10245__A2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09284_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[8\]
+ net678 net674 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08235_ net878 net872 net857 vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__and3_4
XANTENNA_fanout1151_A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout507_A _07452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1249_A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08166_ net903 net966 _04239_ net895 vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_43_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08097_ net1028 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__and2b_1
XFILLER_0_113_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08610__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12405__C _03659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload90 clknet_leaf_52_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload90/Y sky130_fd_sc_hd__clkinv_8
XANTENNA_fanout497_X net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout876_A net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout664_X net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08999_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[14\]
+ net685 net673 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__a22o_1
XANTENNA__09714__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_188_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_188_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13009__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10222__A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09323__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_117_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_117_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_98_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10961_ _06800_ _06801_ _06870_ vssd1 vssd1 vccd1 vccd1 _06946_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout831_X net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12848__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08677__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout929_X net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12700_ net235 net2392 net497 vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__mux2_1
X_13680_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[10\]
+ net286 net384 vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10892_ _06775_ _06886_ _06887_ _04170_ vssd1 vssd1 vccd1 vccd1 _06889_ sky130_fd_sc_hd__a31o_1
XFILLER_0_85_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12631_ net1760 _03663_ _03682_ vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15350_ net1096 vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12562_ net1781 _07812_ _03678_ vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18361__1346 vssd1 vssd1 vccd1 vccd1 _18361__1346/HI net1346 sky130_fd_sc_hd__conb_1
XANTENNA__08105__A_N net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14301_ _04491_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__nor2_1
X_11513_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[23\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[23\]
+ net1032 vssd1 vssd1 vccd1 vccd1 _07424_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13679__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12583__S _03680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15281_ net1192 vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__inv_2
X_12493_ net1675 _07812_ _03673_ vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17020_ clknet_leaf_158_wb_clk_i _02650_ _00716_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_14232_ net1496 _04027_ vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__xor2_1
X_11444_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[30\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[30\]
+ net1033 vssd1 vssd1 vccd1 vccd1 _07356_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_117_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11197__B1 _07129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14163_ _03989_ net907 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[12\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_169_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11375_ net731 _07087_ _07311_ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_169_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09608__D net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13114_ net278 net2510 net448 vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__mux2_1
X_10326_ _05929_ _05983_ _05986_ vssd1 vssd1 vccd1 vccd1 _06347_ sky130_fd_sc_hd__or3_1
X_14094_ _03944_ _03946_ _03959_ vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__o21a_1
X_17922_ clknet_leaf_43_wb_clk_i _03261_ _01618_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13045_ net270 net2468 net456 vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__mux2_1
X_10257_ net1020 _04633_ _04635_ net552 vssd1 vssd1 vccd1 vccd1 _06281_ sky130_fd_sc_hd__a211o_1
XFILLER_0_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1220 net1241 vssd1 vssd1 vccd1 vccd1 net1220 sky130_fd_sc_hd__buf_2
XFILLER_0_56_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1231 net1234 vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__buf_2
X_17853_ clknet_leaf_101_wb_clk_i _03196_ _01549_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[35\]
+ sky130_fd_sc_hd__dfrtp_1
X_10188_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[29\] net903 net965
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[29\] vssd1 vssd1
+ vccd1 vccd1 _06215_ sky130_fd_sc_hd__a22oi_4
Xfanout1242 net1243 vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__buf_4
Xfanout1253 net1255 vssd1 vssd1 vccd1 vccd1 net1253 sky130_fd_sc_hd__buf_4
Xfanout1264 net1279 vssd1 vssd1 vccd1 vccd1 net1264 sky130_fd_sc_hd__clkbuf_2
Xfanout1275 net1276 vssd1 vssd1 vccd1 vccd1 net1275 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_4_14__f_wb_clk_i_X clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16804_ clknet_leaf_181_wb_clk_i _02434_ _00500_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1286 net1287 vssd1 vssd1 vccd1 vccd1 net1286 sky130_fd_sc_hd__clkbuf_4
Xfanout1297 net1298 vssd1 vssd1 vccd1 vccd1 net1297 sky130_fd_sc_hd__buf_4
X_17784_ clknet_leaf_94_wb_clk_i _03127_ _01480_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14996_ net1073 vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__inv_2
XANTENNA__09314__B1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13947_ net910 _03820_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[2\]
+ sky130_fd_sc_hd__nor2_1
X_16735_ clknet_leaf_154_wb_clk_i _02365_ _00431_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09865__A1 _05888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08668__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12758__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09640__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16666_ clknet_leaf_10_wb_clk_i _02296_ _00362_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13878_ net1556 net983 _03775_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[10\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15617_ net1157 vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__inv_2
X_18405_ net1374 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__buf_2
XFILLER_0_146_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12829_ net197 net2853 net481 vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16597_ clknet_leaf_23_wb_clk_i _02227_ _00293_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_173_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18336_ net1325 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XANTENNA__12621__A0 _03646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15548_ net1176 vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09093__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13589__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18267_ clknet_leaf_36_wb_clk_i _03496_ _01962_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_127_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15479_ net1167 vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__inv_2
XANTENNA__12493__S _03673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12346__X _03641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08840__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17218_ clknet_leaf_5_wb_clk_i _02848_ _00914_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18198_ clknet_leaf_36_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[19\]
+ _01893_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08272__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[14\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11188__B1 _07126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold703 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[5\] vssd1
+ vssd1 vccd1 vccd1 net2117 sky130_fd_sc_hd__dlygate4sd3_1
Xhold714 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2128 sky130_fd_sc_hd__dlygate4sd3_1
X_17149_ clknet_leaf_111_wb_clk_i _02779_ _00845_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10307__A _06328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold725 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 net2150 sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net2161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2172 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09971_ _04428_ _05999_ vssd1 vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__xnor2_1
Xhold769 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2183 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08922_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[16\]
+ net676 net625 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[16\]
+ _04976_ vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__a221o_1
XFILLER_0_110_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09553__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08853_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[18\]
+ net590 _04915_ _04920_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[18\]
+ sky130_fd_sc_hd__o22a_4
Xhold1403 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2817 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1414 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 net2828 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1425 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 net2839 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1436 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net2850 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1447 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2861 sky130_fd_sc_hd__dlygate4sd3_1
X_08784_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[19\]
+ net664 net636 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1458 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2872 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1469 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 net2883 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_140_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08659__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08513__D1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout457_A _03712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09405_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[6\]
+ net823 net783 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[6\]
+ _05446_ vssd1 vssd1 vccd1 vccd1 _05449_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_49_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11144__Y _07110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout245_X net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09336_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[7\]
+ net713 net642 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__a22o_1
XANTENNA__09084__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13499__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09267_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[9\]
+ net851 net754 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[9\]
+ _05316_ vssd1 vssd1 vccd1 vccd1 _05317_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout412_X net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08831__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08218_ net881 net866 _04294_ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__and3_4
XFILLER_0_90_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09198_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[10\]
+ net690 net676 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[10\]
+ _05250_ vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__a221o_1
XANTENNA__11179__B1 _07127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09709__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08149_ net1022 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[5\]
+ _04231_ vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__nor3_2
XTAP_TAPCELL_ROW_75_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11708__D_N team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_892 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11160_ _07039_ _07081_ vssd1 vssd1 vccd1 vccd1 _07126_ sky130_fd_sc_hd__nor2_4
Xclkload190 clknet_leaf_99_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload190/Y sky130_fd_sc_hd__inv_6
XANTENNA_fanout781_X net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10111_ _06135_ _06138_ net513 vssd1 vssd1 vccd1 vccd1 _06139_ sky130_fd_sc_hd__mux2_1
X_11091_ _04161_ _07056_ _07057_ _07053_ vssd1 vssd1 vccd1 vccd1 _07058_ sky130_fd_sc_hd__a31o_2
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10651__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_164_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09544__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10042_ net520 _06070_ vssd1 vssd1 vccd1 vccd1 _06071_ sky130_fd_sc_hd__nand2_1
Xhold30 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[16\]
+ vssd1 vssd1 vccd1 vccd1 net1444 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08898__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold41 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[11\] vssd1 vssd1
+ vccd1 vccd1 net1455 sky130_fd_sc_hd__dlygate4sd3_1
X_14850_ net1193 vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__inv_2
Xhold52 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[8\]
+ vssd1 vssd1 vccd1 vccd1 net1466 sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[15\]
+ vssd1 vssd1 vccd1 vccd1 net1477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[12\]
+ vssd1 vssd1 vccd1 vccd1 net1488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[16\]
+ vssd1 vssd1 vccd1 vccd1 net1499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[22\]
+ vssd1 vssd1 vccd1 vccd1 net1510 sky130_fd_sc_hd__dlygate4sd3_1
X_13801_ net1560 net975 net724 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[12\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_98_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11990__B _07798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input18_A DAT_I[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14781_ net1089 vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__inv_2
X_11993_ _07716_ _07787_ _07804_ vssd1 vssd1 vccd1 vccd1 _07805_ sky130_fd_sc_hd__and3_1
XANTENNA__11482__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16520_ clknet_leaf_204_wb_clk_i _02150_ _00216_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13732_ net921 _06756_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[0\]
+ sky130_fd_sc_hd__nor2_1
X_10944_ _06875_ _06931_ net1043 vssd1 vssd1 vccd1 vccd1 _06932_ sky130_fd_sc_hd__and3b_1
X_16451_ clknet_leaf_199_wb_clk_i _02081_ _00147_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13663_ net2449 net222 net385 vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__mux2_1
X_10875_ _06801_ _06871_ vssd1 vssd1 vccd1 vccd1 _06872_ sky130_fd_sc_hd__or2_1
X_15402_ net1131 vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__inv_2
X_12614_ _03661_ net1814 net201 vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16382_ clknet_leaf_163_wb_clk_i _02012_ _00078_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13594_ net2656 net195 net394 vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__mux2_1
XANTENNA__09075__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_85_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_18121_ clknet_leaf_45_wb_clk_i _00035_ _01817_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_15333_ net1203 vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13710__B _06591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12545_ _07857_ net2066 net207 vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08822__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13202__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_18052_ net1037 _03390_ _01748_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15264_ net1105 vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__inv_2
X_12476_ net1745 net500 net210 vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__mux2_1
X_17003_ clknet_leaf_185_wb_clk_i _02633_ _00699_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_14215_ _04013_ net728 _04012_ vssd1 vssd1 vccd1 vccd1 _00009_ sky130_fd_sc_hd__and3b_1
X_11427_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[1\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[0\]
+ vssd1 vssd1 vccd1 vccd1 _07342_ sky130_fd_sc_hd__or2_1
XANTENNA_5 _07434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15195_ net1100 vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14146_ team_05_WB.instance_to_wrap.CPU_DAT_O\[29\] net504 net912 vssd1 vssd1 vccd1
+ vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[29\] sky130_fd_sc_hd__and3_1
X_11358_ _07289_ _07293_ _07298_ _07299_ vssd1 vssd1 vccd1 vccd1 _07300_ sky130_fd_sc_hd__a211o_1
XFILLER_0_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10309_ net531 _06230_ _06330_ vssd1 vssd1 vccd1 vccd1 _06331_ sky130_fd_sc_hd__a21o_1
X_14077_ _03943_ _03944_ vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__or2_1
X_11289_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[121\] _07099_
+ _07123_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[97\] vssd1 vssd1
+ vccd1 vccd1 _07249_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_5_Left_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09535__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17905_ clknet_leaf_100_wb_clk_i _03248_ _01601_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13028_ _04253_ net562 _03708_ vssd1 vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__or3_4
XANTENNA__08889__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1050 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read vssd1
+ vssd1 vccd1 vccd1 net1050 sky130_fd_sc_hd__clkbuf_4
Xfanout1061 net1064 vssd1 vssd1 vccd1 vccd1 net1061 sky130_fd_sc_hd__buf_2
X_17836_ clknet_leaf_77_wb_clk_i _03179_ _01532_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[82\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1072 net1108 vssd1 vssd1 vccd1 vccd1 net1072 sky130_fd_sc_hd__clkbuf_4
Xfanout1083 net1086 vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__buf_4
Xfanout1094 net1107 vssd1 vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17767_ clknet_leaf_87_wb_clk_i _03110_ _01463_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12488__S _03674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09299__C1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14979_ net1203 vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16718_ clknet_leaf_175_wb_clk_i _02348_ _00414_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17698_ clknet_leaf_95_wb_clk_i _03041_ _01394_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[72\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08267__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[26\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16649_ clknet_leaf_19_wb_clk_i _02279_ _00345_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13460__X _03728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09121_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[12\]
+ net778 net760 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[12\]
+ _05176_ vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_44_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18319_ net1411 vssd1 vssd1 vccd1 vccd1 gpio_oeb[34] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_44_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08813__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13112__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09052_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[13\]
+ net710 net698 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[13\]
+ _05110_ vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_96_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12951__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold500 net111 vssd1 vssd1 vccd1 vccd1 net1914 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold511 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1925 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout205_A net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold522 team_05_WB.instance_to_wrap.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 net1936
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold533 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 net1947 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold544 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net1958 sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net1969 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10384__B2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[21\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold566 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net1980 sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net1991 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold588 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 net2002 sky130_fd_sc_hd__dlygate4sd3_1
X_09954_ _05980_ _05981_ vssd1 vssd1 vccd1 vccd1 _05983_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10324__X _06346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold599 _03301_ vssd1 vssd1 vccd1 vccd1 net2013 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14170__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09526__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08905_ _04967_ _04969_ vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__nor2_4
XANTENNA__11139__Y _07105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09885_ _04553_ _04533_ vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout574_A net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1200 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2614 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1211 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net2625 sky130_fd_sc_hd__dlygate4sd3_1
X_18360__1345 vssd1 vssd1 vccd1 vccd1 _18360__1345/HI net1345 sky130_fd_sc_hd__conb_1
Xhold1222 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2636 sky130_fd_sc_hd__dlygate4sd3_1
X_08836_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[18\]
+ net777 net770 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[18\]
+ _04903_ vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__a221o_1
Xhold1233 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2647 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1244 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net2658 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1255 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2669 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1266 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 net2680 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13086__A0 _06655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12398__S _07852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08767_ _04344_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[21\]
+ _04362_ vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__o21ai_1
Xhold1277 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2691 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14179__A team_05_WB.instance_to_wrap.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold1288 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2702 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout741_A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1299 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2713 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout839_A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_68_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08698_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[22\]
+ net689 net654 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_68_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09711__D net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout627_X net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14907__A net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10660_ net529 _06595_ _06064_ vssd1 vssd1 vccd1 vccd1 _06664_ sky130_fd_sc_hd__o21a_1
XFILLER_0_153_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09319_ _05360_ _05363_ _05365_ _05366_ vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__or4_1
XFILLER_0_165_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12061__A1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[11\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10591_ _05285_ net511 _06284_ _06510_ vssd1 vssd1 vccd1 vccd1 _06599_ sky130_fd_sc_hd__o22a_1
XFILLER_0_51_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13022__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12330_ _03615_ _03618_ _03624_ _03610_ vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__or4b_1
XFILLER_0_145_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13010__A0 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12261_ _07947_ _07959_ _03553_ vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14000_ _03867_ _03870_ vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__nand2_1
X_11212_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[13\] _07105_
+ _07169_ _07175_ vssd1 vssd1 vccd1 vccd1 _07176_ sky130_fd_sc_hd__a211o_1
XANTENNA__09765__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12192_ _07987_ _07995_ _07998_ _08001_ _08002_ vssd1 vssd1 vccd1 vccd1 _08004_ sky130_fd_sc_hd__a32o_1
XANTENNA__10375__A1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10375__B2 _06355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11143_ _07039_ _07083_ vssd1 vssd1 vccd1 vccd1 _07109_ sky130_fd_sc_hd__nor2_4
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 ADR_O[0] sky130_fd_sc_hd__clkbuf_4
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 ADR_O[1] sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_132_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_132_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__clkbuf_4
X_11074_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[2\] team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[0\]
+ _07033_ vssd1 vssd1 vccd1 vccd1 _07041_ sky130_fd_sc_hd__a21oi_1
X_15951_ net1302 vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__inv_2
X_10025_ net1018 _05923_ vssd1 vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__nor2_1
X_14902_ net1091 vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__inv_2
X_15882_ net1290 vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17621_ clknet_leaf_59_wb_clk_i _02992_ _01317_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14833_ net1188 vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17552_ clknet_leaf_58_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[23\]
+ _01248_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14764_ net1109 vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__inv_2
XANTENNA__10410__A net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11976_ net501 _07718_ vssd1 vssd1 vccd1 vccd1 _07788_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11627__B2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09296__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13715_ net899 _06500_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[15\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_38_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16503_ clknet_leaf_143_wb_clk_i _02133_ _00199_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10927_ _05906_ _06917_ vssd1 vssd1 vccd1 vccd1 _06918_ sky130_fd_sc_hd__or2_4
X_17483_ clknet_leaf_37_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[18\]
+ _01179_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14695_ net1104 vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13721__A _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13646_ net2429 net292 net388 vssd1 vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__mux2_1
X_16434_ clknet_leaf_136_wb_clk_i _02064_ _00130_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10858_ _06826_ _06854_ vssd1 vssd1 vccd1 vccd1 _06855_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09048__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08256__B1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16365_ clknet_leaf_159_wb_clk_i _01995_ _00061_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13577_ net2726 net276 net399 vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__mux2_1
X_10789_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[25\] net1040 vssd1
+ vssd1 vccd1 vccd1 _06786_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18104_ clknet_leaf_52_wb_clk_i _03427_ _01800_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[21\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_143_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15316_ net1067 vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__inv_2
X_12528_ _03663_ net1829 _03675_ vssd1 vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__mux2_1
X_16296_ net1147 vssd1 vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18035_ clknet_leaf_97_wb_clk_i _03374_ _01731_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_15247_ net1281 vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__inv_2
X_12459_ net1710 _03663_ _03670_ vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__mux2_1
XANTENNA__12771__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09756__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire375_A _05397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15178_ net1122 vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09220__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11563__B1 _07394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14129_ net1577 net507 _03991_ vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_123_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout309 net312 vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09508__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11315__B1 _07124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_77_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09670_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[1\]
+ net876 net867 net860 vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__and4_1
XFILLER_0_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08621_ _04682_ _04693_ _04694_ _04695_ vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__or4_1
X_17819_ clknet_leaf_76_wb_clk_i _03162_ _01515_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[65\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13107__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08552_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[26\]
+ net831 _04628_ net856 vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__a211o_1
XANTENNA__10320__A net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11618__B2 _07478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09287__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_59_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12946__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08483_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[27\]
+ net705 net641 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[27\]
+ _04557_ vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__a221o_1
XANTENNA__14727__A net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08284__X _04366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12043__A1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[23\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08247__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10466__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout322_A net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1064_A net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09104_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[12\]
+ net664 net636 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09035_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[14\]
+ net834 net734 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1231_A net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout208_X net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_68_Left_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold330 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[126\] vssd1 vssd1
+ vccd1 vccd1 net1744 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold341 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[17\] vssd1 vssd1
+ vccd1 vccd1 net1755 sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[14\] vssd1 vssd1
+ vccd1 vccd1 net1766 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09211__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout691_A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold363 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[16\] vssd1 vssd1
+ vccd1 vccd1 net1777 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout789_A _04400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold374 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[96\] vssd1 vssd1
+ vccd1 vccd1 net1788 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold385 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[38\] vssd1 vssd1
+ vccd1 vccd1 net1799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[107\] vssd1 vssd1
+ vccd1 vccd1 net1810 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout810 net813 vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09706__D net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout821 _04387_ vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__clkbuf_8
X_09937_ _05831_ _05962_ _05965_ _05832_ vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__o211ai_1
Xfanout832 _04382_ vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__buf_4
Xfanout843 net844 vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__buf_4
XANTENNA__11306__B1 _07265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout577_X net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout956_A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout854 _04367_ vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__clkbuf_4
Xfanout865 net866 vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout876 net882 vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__clkbuf_2
X_09868_ _05895_ _05896_ vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__or2_1
Xfanout887 _04281_ vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__buf_1
Xfanout898 _04248_ vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__buf_2
Xhold1030 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1041 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net2455 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1052 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 net2466 sky130_fd_sc_hd__dlygate4sd3_1
X_08819_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[18\]
+ net711 net629 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[18\]
+ _04887_ vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__a221o_1
Xhold1063 net105 vssd1 vssd1 vccd1 vccd1 net2477 sky130_fd_sc_hd__dlygate4sd3_1
X_09799_ _05144_ _05123_ vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__and2b_1
Xhold1074 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2488 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout744_X net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09722__C net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1085 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net2499 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13017__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1096 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2510 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12806__A0 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_77_Left_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ _07639_ _07640_ _07629_ vssd1 vssd1 vccd1 vccd1 _07642_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_29_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09278__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08486__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11761_ _07569_ _07571_ vssd1 vssd1 vccd1 vccd1 _07573_ sky130_fd_sc_hd__nand2_1
XANTENNA__12856__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13500_ net2050 net239 net406 vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__mux2_1
XANTENNA__10293__B1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10712_ _05806_ _06054_ vssd1 vssd1 vccd1 vccd1 _06713_ sky130_fd_sc_hd__nand2_1
X_14480_ net1182 vssd1 vssd1 vccd1 vccd1 _00110_ sky130_fd_sc_hd__inv_2
X_11692_ net73 net71 net74 _07504_ vssd1 vssd1 vccd1 vccd1 _07505_ sky130_fd_sc_hd__and4_1
X_13431_ net2550 net220 net414 vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__mux2_1
X_10643_ net524 _06581_ _06647_ vssd1 vssd1 vccd1 vccd1 _06648_ sky130_fd_sc_hd__a21o_1
XFILLER_0_165_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16150_ net1263 vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13362_ net2224 net198 net421 vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_172_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10574_ _06431_ net332 _06582_ net335 _06579_ vssd1 vssd1 vccd1 vccd1 _06583_ sky130_fd_sc_hd__o221a_1
XANTENNA__09450__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10596__B2 _06603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15101_ net1089 vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__inv_2
X_12313_ net250 net251 _03602_ vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13687__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16081_ net1259 vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__inv_2
XANTENNA__12591__S net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_86_Left_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13293_ net324 net2075 net432 vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__mux2_1
XANTENNA__09737__Y team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15032_ net1242 vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__inv_2
XANTENNA__09738__B1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12244_ _03524_ _03527_ _03518_ vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09466__A net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_111_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12175_ _07941_ _07986_ vssd1 vssd1 vccd1 vccd1 _07987_ sky130_fd_sc_hd__xor2_1
XANTENNA__10405__A net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11000__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09616__D net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11126_ _07038_ _07068_ _07073_ vssd1 vssd1 vccd1 vccd1 _07092_ sky130_fd_sc_hd__and3_4
X_16983_ clknet_leaf_143_wb_clk_i _02613_ _00679_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10124__B net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13716__A _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09472__Y team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11057_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[7\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[6\]
+ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[9\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[8\]
+ vssd1 vssd1 vccd1 vccd1 _07024_ sky130_fd_sc_hd__or4_1
X_15934_ net1272 vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__inv_2
XANTENNA__09913__B net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_95_Left_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10008_ _04944_ net364 vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__or2_1
X_15865_ net1270 vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__inv_2
X_17604_ clknet_leaf_80_wb_clk_i _02975_ _01300_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14816_ net1198 vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__inv_2
XANTENNA__10140__A net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15796_ net1300 vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__inv_2
XANTENNA__09269__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17535_ clknet_leaf_79_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[6\]
+ _01231_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11959_ _07767_ _07769_ _07765_ vssd1 vssd1 vccd1 vccd1 _07771_ sky130_fd_sc_hd__o21a_1
XANTENNA__08477__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14747_ net1095 vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__inv_2
XANTENNA__12766__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11523__X _07434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17466_ clknet_leaf_39_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[1\]
+ _01162_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14678_ net1085 vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12025__A1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[19\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16417_ clknet_leaf_149_wb_clk_i _02047_ _00113_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13629_ net2596 net220 net391 vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17397_ clknet_leaf_60_wb_clk_i net1430 _01093_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08264__B team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[22\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_150_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16348_ clknet_leaf_154_wb_clk_i _01978_ _00044_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13597__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16279_ net1155 vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__inv_2
XANTENNA__14282__A _06572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13525__A1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18018_ clknet_leaf_96_wb_clk_i _03357_ _01714_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_130_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09376__A net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire378_X net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08280__A net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08401__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09722_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[0\]
+ net1017 net950 net929 vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__and4_1
X_09653_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[1\]
+ net849 net795 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_87_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08604_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[24\]
+ net653 net595 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__a22o_1
X_09584_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[2\]
+ net1015 net941 net932 vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__and4_1
XFILLER_0_167_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08535_ _04597_ _04598_ _04600_ _04611_ vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__or4_2
XFILLER_0_77_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08468__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout537_A net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1181_A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11433__X _07346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1279_A net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08466_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[28\]
+ net839 net735 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11152__Y _07118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13213__A0 _06570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout704_A _04292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08397_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[29\]
+ net633 net611 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[29\]
+ _04472_ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__a221o_1
XFILLER_0_162_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10578__A1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09432__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10578__B2 _04175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1234_X net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08902__B _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13300__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09018_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[14\] _04354_
+ vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10290_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[24\] _06099_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[25\]
+ vssd1 vssd1 vccd1 vccd1 _06313_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08190__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout694_X net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09717__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold160 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[30\]
+ vssd1 vssd1 vccd1 vccd1 net1574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[7\] vssd1 vssd1
+ vccd1 vccd1 net1585 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold182 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[14\]
+ vssd1 vssd1 vccd1 vccd1 net1596 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold193 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[22\]
+ vssd1 vssd1 vccd1 vccd1 net1607 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout861_X net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout959_X net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout640 net643 vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_109_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout651 _04309_ vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout662 net663 vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__clkbuf_8
X_13980_ _03828_ _03831_ _03851_ vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__o21ba_1
XANTENNA__11982__C _07793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout673 net675 vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09499__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout684 net685 vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__clkbuf_8
Xfanout695 net698 vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__clkbuf_8
X_12931_ net194 net2806 net469 vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_126_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15650_ net1250 vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__inv_2
X_12862_ net197 net2867 net477 vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__mux2_1
X_14601_ net1215 vssd1 vssd1 vccd1 vccd1 _00231_ sky130_fd_sc_hd__inv_2
X_11813_ _07620_ _07623_ _07624_ vssd1 vssd1 vccd1 vccd1 _07625_ sky130_fd_sc_hd__or3_2
X_15581_ net1250 vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08459__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12439__X _03670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12586__S _03680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[10\] _04255_
+ vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__nor2_1
XANTENNA__14367__A _04094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17320_ clknet_leaf_1_wb_clk_i _02950_ _01016_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_14532_ net1208 vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_174_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _07533_ _07546_ vssd1 vssd1 vccd1 vccd1 _07556_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_174_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13204__A0 _06404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14463_ net1178 vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__inv_2
X_17251_ clknet_leaf_199_wb_clk_i _02881_ _00947_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11675_ _07489_ vssd1 vssd1 vccd1 vccd1 _07490_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_12_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_1112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13414_ net2008 net278 net416 vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16202_ net1077 vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__inv_2
X_10626_ net1020 _05375_ _05377_ net551 vssd1 vssd1 vccd1 vccd1 _06632_ sky130_fd_sc_hd__a211o_1
X_17182_ clknet_leaf_184_wb_clk_i _02812_ _00878_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14394_ net1508 vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10569__A1 _05208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14373__Y _04146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09423__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16133_ net1292 vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13345_ net270 net2776 net424 vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__mux2_1
XANTENNA__15198__A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11230__A2 _07123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10557_ _06565_ _06566_ net536 vssd1 vssd1 vccd1 vccd1 _06567_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08812__B net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13210__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16064_ net1259 vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__inv_2
X_13276_ net266 net2448 net432 vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__mux2_1
X_10488_ _05935_ _05964_ vssd1 vssd1 vccd1 vccd1 _06501_ sky130_fd_sc_hd__xor2_1
X_15015_ net1242 vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__inv_2
X_12227_ _08012_ _08016_ _08017_ vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__and3_1
XANTENNA__14830__A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12158_ _07969_ vssd1 vssd1 vccd1 vccd1 _07970_ sky130_fd_sc_hd__inv_2
XANTENNA__17914__Q team_05_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17563__D team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11109_ _07073_ _07075_ vssd1 vssd1 vccd1 vccd1 _07076_ sky130_fd_sc_hd__nand2_2
XFILLER_0_75_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16966_ clknet_leaf_116_wb_clk_i _02596_ _00662_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12089_ _07898_ _07900_ vssd1 vssd1 vccd1 vccd1 _07901_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_34_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15917_ net1288 vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__inv_2
XANTENNA__11297__A2 _07109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12494__A1 _03663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08698__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16897_ clknet_leaf_147_wb_clk_i _02527_ _00593_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15848_ net1275 vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11049__A2 _06706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12496__S _03674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15779_ net1305 vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__inv_2
XANTENNA__12349__X _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08320_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[31\]
+ net788 net783 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__a22o_1
X_17518_ clknet_leaf_74_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[21\]
+ _01214_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_115_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09662__A2 _04366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12509__B _03659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08251_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[31\]
+ net692 net618 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[31\]
+ _04333_ vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__a221o_1
XFILLER_0_89_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17449_ clknet_leaf_47_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[17\]
+ _01145_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08870__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08182_ _04258_ _04263_ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__nand2_4
XANTENNA__09414__A2 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11221__A2 _07097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13120__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10316__Y _06338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10045__A _04573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10732__A1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout487_A _03703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10732__B2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09705_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[0\]
+ net591 vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__nor2_1
XANTENNA__11147__Y _07113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11288__A2 _07111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12485__A1 _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08689__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout654_A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08169__B team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09636_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[13\] net968
+ _04268_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[8\] _05670_
+ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[1\]
+ sky130_fd_sc_hd__a221o_2
XTAP_TAPCELL_ROW_104_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09567_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[2\]
+ net947 net939 net930 vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout821_A _04387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout442_X net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11163__X _07129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08518_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[26\]
+ net693 net623 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__a22o_1
X_09498_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[4\]
+ net705 net653 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__a22o_1
XANTENNA__09653__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08449_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[28\]
+ net631 net627 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[28\]
+ _04527_ vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_863 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08861__B1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout707_X net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11460_ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[6\] _07370_ net1002
+ vssd1 vssd1 vccd1 vccd1 _07371_ sky130_fd_sc_hd__mux2_2
XFILLER_0_18_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09405__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10411_ _06425_ _06427_ net556 vssd1 vssd1 vccd1 vccd1 _06428_ sky130_fd_sc_hd__a21o_1
XANTENNA__11212__A2 _07105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11391_ _04165_ _07321_ vssd1 vssd1 vccd1 vccd1 _07322_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08613__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13030__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10420__B1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13130_ net191 net2880 net446 vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__mux2_1
X_10342_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[23\] _06098_ vssd1
+ vssd1 vccd1 vccd1 _06363_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_78_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13061_ _04257_ _04261_ net562 vssd1 vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__or3_4
X_10273_ _05905_ _06295_ vssd1 vssd1 vccd1 vccd1 _06296_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12012_ net343 _07758_ _07772_ _07823_ vssd1 vssd1 vccd1 vccd1 _07824_ sky130_fd_sc_hd__a31o_1
XANTENNA_input48_A wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11485__S net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_39_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08392__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16820_ clknet_leaf_115_wb_clk_i _02450_ _00516_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10242__X _06267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout470 net471 vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__buf_4
Xfanout481 net482 vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_6_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11279__A2 _07119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12476__A1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16751_ clknet_leaf_134_wb_clk_i _02381_ _00447_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout492 net493 vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__buf_6
X_13963_ _03834_ _03835_ _03805_ vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15702_ net1153 vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__inv_2
X_12914_ net280 net2294 net472 vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__mux2_1
X_13894_ net1598 net981 _03783_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[18\]
+ sky130_fd_sc_hd__o21a_1
X_16682_ clknet_leaf_196_wb_clk_i _02312_ _00378_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13713__B _06540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12845_ net271 net2907 net480 vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__mux2_1
X_15633_ net1245 vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09629__C1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08366__Y _04447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13205__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18352_ net1337 vssd1 vssd1 vccd1 vccd1 la_data_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_57_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12776_ net269 net2508 net488 vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__mux2_1
X_15564_ net1246 vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_14_Left_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17303_ clknet_leaf_146_wb_clk_i _02933_ _00999_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11727_ _07479_ _07538_ _07537_ _07530_ _07519_ vssd1 vssd1 vccd1 vccd1 _07539_ sky130_fd_sc_hd__o2111a_1
X_14515_ net1215 vssd1 vssd1 vccd1 vccd1 _00145_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_3_0_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18283_ net107 vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__clkbuf_1
X_15495_ net1159 vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14825__A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_868 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17234_ clknet_leaf_133_wb_clk_i _02864_ _00930_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11658_ net4 net990 net917 net1687 vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__o22a_1
X_14446_ net1189 vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10609_ _05818_ _06615_ _05819_ net511 vssd1 vssd1 vccd1 vccd1 _06616_ sky130_fd_sc_hd__o2bb2a_1
X_14377_ net1536 vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12400__A1 _03650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11203__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17165_ clknet_leaf_161_wb_clk_i _02795_ _00861_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08604__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09638__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11589_ team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.state\[1\] team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.state\[0\]
+ net1048 team_05_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 _07470_ sky130_fd_sc_hd__and4b_4
XFILLER_0_141_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold907 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net2321 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16116_ net1134 vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__inv_2
XANTENNA__10411__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold918 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2332 sky130_fd_sc_hd__dlygate4sd3_1
X_13328_ team_05_WB.instance_to_wrap.total_design.core.instr_fetch _04258_ _04261_
+ _03702_ vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__or4_4
XFILLER_0_122_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17096_ clknet_leaf_197_wb_clk_i _02726_ _00792_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold929 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 net2343 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16047_ net1287 vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__inv_2
X_13259_ net321 net2065 net436 vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_23_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10714__A1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08383__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17998_ clknet_leaf_82_wb_clk_i _03337_ _01694_ vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12467__A1 _07821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16949_ clknet_leaf_116_wb_clk_i _02579_ _00645_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_84_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10478__A0 _06338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09421_ _05442_ _05463_ vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13115__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09352_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[19\] net967
+ _05398_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[27\] vssd1
+ vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__a22oi_1
XANTENNA__09096__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08303_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[31\]
+ net827 net823 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09283_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[8\]
+ net689 net604 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__a22o_1
XANTENNA__08843__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12954__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout235_A net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11550__B_N _07409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10650__B1 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08234_ net880 net875 _04287_ vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__and3_1
XFILLER_0_173_974 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08165_ net962 net955 vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout402_A net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08096_ net1029 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[13\]
+ net976 _04197_ vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload80 clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload80/Y sky130_fd_sc_hd__inv_8
XFILLER_0_101_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload91 clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload91/Y sky130_fd_sc_hd__inv_12
XANTENNA__15566__A net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1311_A net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10166__C1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout771_A _04406_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout392_X net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08374__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout869_A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08998_ _05058_ vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__inv_2
XANTENNA__09714__D net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12458__A1 _07812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09859__C1 _05887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout657_X net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10222__B _06247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_170_Right_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10960_ _06800_ _06801_ _06870_ vssd1 vssd1 vccd1 vccd1 _06945_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09619_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[2\]
+ net695 _05638_ _05643_ _05653_ vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__a2111o_1
X_10891_ _06775_ _06886_ _06887_ vssd1 vssd1 vccd1 vccd1 _06888_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout824_X net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13025__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12630_ net1691 _07812_ _03682_ vssd1 vssd1 vccd1 vccd1 _03015_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_157_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_157_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09626__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12561_ _03645_ net1886 net207 vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12630__A1 _07812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12864__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11512_ _07348_ _07353_ _07422_ vssd1 vssd1 vccd1 vccd1 _07423_ sky130_fd_sc_hd__or3_1
X_14300_ net380 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__nor2_1
X_15280_ net1183 vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__inv_2
X_12492_ net1704 _03645_ net210 vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14231_ team_05_WB.instance_to_wrap.total_design.keypad0.counter\[16\] team_05_WB.instance_to_wrap.total_design.keypad0.counter\[17\]
+ _04026_ vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__and3_1
XFILLER_0_108_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11443_ net1928 net1004 _07348_ net727 vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14162_ _03980_ net907 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[11\]
+ sky130_fd_sc_hd__nor2_1
X_11374_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[5\] net732
+ vssd1 vssd1 vccd1 vccd1 _07311_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_169_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_169_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13113_ net282 net2155 net449 vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__mux2_1
X_10325_ net2103 net235 net540 vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__mux2_1
X_14093_ _03944_ _03946_ _03959_ vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__or3_1
X_17921_ clknet_leaf_35_wb_clk_i _03260_ _01617_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13044_ net269 net2599 net456 vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__mux2_1
X_10256_ _06139_ _06148_ net530 vssd1 vssd1 vccd1 vccd1 _06280_ sky130_fd_sc_hd__mux2_1
XANTENNA__13708__B _06623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1210 net1211 vssd1 vssd1 vccd1 vccd1 net1210 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09562__A1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[14\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1221 net1222 vssd1 vssd1 vccd1 vccd1 net1221 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17852_ clknet_leaf_88_wb_clk_i _03195_ _01548_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09562__B2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[22\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1232 net1234 vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__buf_4
X_10187_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[29\] _06102_ vssd1
+ vssd1 vccd1 vccd1 _06214_ sky130_fd_sc_hd__xnor2_2
Xfanout1243 net1312 vssd1 vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__clkbuf_4
Xfanout1254 net1255 vssd1 vssd1 vccd1 vccd1 net1254 sky130_fd_sc_hd__clkbuf_2
Xfanout1265 net1268 vssd1 vssd1 vccd1 vccd1 net1265 sky130_fd_sc_hd__buf_4
X_16803_ clknet_leaf_198_wb_clk_i _02433_ _00499_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1276 net1278 vssd1 vssd1 vccd1 vccd1 net1276 sky130_fd_sc_hd__buf_4
XANTENNA__12449__A1 _03646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17783_ clknet_leaf_84_wb_clk_i _03126_ _01479_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1287 net1312 vssd1 vssd1 vccd1 vccd1 net1287 sky130_fd_sc_hd__buf_4
X_14995_ net1217 vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__inv_2
Xfanout1298 net1311 vssd1 vssd1 vccd1 vccd1 net1298 sky130_fd_sc_hd__buf_2
XANTENNA__13724__A net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16734_ clknet_leaf_184_wb_clk_i _02364_ _00430_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13946_ net1937 net507 _03819_ vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09640__C net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16665_ clknet_leaf_10_wb_clk_i _02295_ _00361_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13877_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[10\]
+ net559 net577 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[10\]
+ net988 vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__a221o_1
X_18404_ net915 vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_1
X_15616_ net1157 vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09078__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12828_ net563 _03695_ _03702_ vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__or3_1
X_16596_ clknet_leaf_128_wb_clk_i _02226_ _00292_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_146_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18335_ net1324 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
X_15547_ net1116 vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__inv_2
XANTENNA__12774__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08825__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12759_ net305 net2266 net493 vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18266_ clknet_leaf_33_wb_clk_i _03495_ _01961_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[20\]
+ sky130_fd_sc_hd__dfrtp_4
X_15478_ net1167 vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14374__A1 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17217_ clknet_leaf_147_wb_clk_i _02847_ _00913_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_14429_ net1091 vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__inv_2
X_18197_ clknet_leaf_36_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[18\]
+ _01892_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17148_ clknet_leaf_157_wb_clk_i _02778_ _00844_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold704 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net2118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold715 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net2129 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09250__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold726 net113 vssd1 vssd1 vccd1 vccd1 net2140 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_31_Left_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold737 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net2151 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09970_ _04471_ _05998_ _05926_ vssd1 vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__o21a_1
Xhold748 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 net2162 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12362__X _03657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17079_ clknet_leaf_146_wb_clk_i _02709_ _00775_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold759 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net2173 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire360_X net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08921_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[16\]
+ net606 _04985_ net719 vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__a211o_1
XANTENNA__09002__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08356__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10699__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08852_ _04904_ _04917_ _04918_ _04919_ vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_51_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1404 team_05_WB.instance_to_wrap.wishbone.curr_state\[2\] vssd1 vssd1 vccd1 vccd1
+ net2818 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1415 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net2829 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1426 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net2840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1437 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2851 sky130_fd_sc_hd__dlygate4sd3_1
X_08783_ _04847_ _04849_ _04851_ _04853_ vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__or4_1
XFILLER_0_137_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1448 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2862 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12949__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08108__A2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1459 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 net2873 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout352_A _03717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09404_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[6\]
+ net830 net772 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[6\]
+ _05447_ vssd1 vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1094_A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14168__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_722 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09069__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11995__A1_N _07474_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09335_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[7\]
+ net674 net615 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[7\]
+ _05380_ vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__a221o_1
XANTENNA__08816__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1261_A net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout617_A net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09266_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[9\]
+ net812 net739 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13800__C net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11160__Y _07126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_950 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08217_ net878 net870 net865 vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__and3_1
XFILLER_0_172_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09197_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[10\]
+ net621 net606 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout405_X net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09709__D net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08148_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[3\] team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[2\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[1\] team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__or4bb_4
XANTENNA__09241__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08595__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08079_ net1027 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__and2b_1
Xclkload180 clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload180/Y sky130_fd_sc_hd__inv_8
Xclkload191 clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload191/Y sky130_fd_sc_hd__inv_8
XFILLER_0_30_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10110_ _06136_ _06137_ vssd1 vssd1 vccd1 vccd1 _06138_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_112_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11090_ _07032_ _07044_ _07055_ vssd1 vssd1 vccd1 vccd1 _07057_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_8_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout774_X net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_164_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_164_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10041_ net380 net367 vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__nor2_1
XANTENNA_hold564_A team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold20 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[4\]
+ vssd1 vssd1 vccd1 vccd1 net1434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[3\]
+ vssd1 vssd1 vccd1 vccd1 net1445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[18\]
+ vssd1 vssd1 vccd1 vccd1 net1456 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[21\] vssd1 vssd1
+ vccd1 vccd1 net1467 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[19\] vssd1 vssd1
+ vccd1 vccd1 net1478 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12859__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold75 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[18\] vssd1 vssd1
+ vccd1 vccd1 net1489 sky130_fd_sc_hd__dlygate4sd3_1
X_13800_ net1566 net976 net725 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[11\]
+ sky130_fd_sc_hd__and3_1
Xhold86 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[12\]
+ vssd1 vssd1 vccd1 vccd1 net1500 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11616__X _07478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold97 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[11\]
+ vssd1 vssd1 vccd1 vccd1 net1511 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11990__C _07797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11992_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[25\] net995 net548
+ vssd1 vssd1 vccd1 vccd1 _07804_ sky130_fd_sc_hd__a21oi_1
X_14780_ net1063 vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__inv_2
X_13731_ net899 _05921_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[31\]
+ sky130_fd_sc_hd__nor2_1
X_10943_ _06793_ _06794_ _06796_ _06874_ vssd1 vssd1 vccd1 vccd1 _06931_ sky130_fd_sc_hd__a211o_1
XFILLER_0_58_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10379__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_28_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_85_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16450_ clknet_leaf_15_wb_clk_i _02080_ _00146_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10874_ _06802_ _06869_ _06800_ vssd1 vssd1 vccd1 vccd1 _06871_ sky130_fd_sc_hd__a21oi_1
X_13662_ net2161 net221 net386 vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15401_ net1222 vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__inv_2
X_12613_ net500 net2095 net201 vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12594__S net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13593_ net2570 net197 net394 vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__mux2_1
X_16381_ clknet_leaf_129_wb_clk_i _02011_ _00077_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18120_ clknet_leaf_46_wb_clk_i _00034_ _01816_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_12544_ _07858_ _07862_ _03659_ vssd1 vssd1 vccd1 vccd1 _03679_ sky130_fd_sc_hd__nand3b_1
XANTENNA__10614__B1 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15332_ net1237 vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09480__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18051_ net1037 _03389_ _01747_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[6\]
+ sky130_fd_sc_hd__dfrtp_2
X_12475_ net919 _07860_ _07863_ _03659_ vssd1 vssd1 vccd1 vccd1 _03674_ sky130_fd_sc_hd__and4b_4
X_15263_ net1179 vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17002_ clknet_leaf_195_wb_clk_i _02632_ _00698_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11426_ _07314_ _07341_ net730 vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__o21bai_1
X_14214_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[12\] _04011_
+ vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__and2_1
X_15194_ net1055 vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_6 team_05_WB.instance_to_wrap.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_54_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_123_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14145_ team_05_WB.instance_to_wrap.CPU_DAT_O\[28\] net504 net912 vssd1 vssd1 vccd1
+ vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[28\] sky130_fd_sc_hd__and3_1
XANTENNA__08586__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11357_ _04216_ _07289_ vssd1 vssd1 vccd1 vccd1 _07299_ sky130_fd_sc_hd__nor2_1
XANTENNA__13719__A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09916__B _05731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08991__C1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10308_ net524 _06239_ net333 vssd1 vssd1 vccd1 vccd1 _06330_ sky130_fd_sc_hd__a21o_1
X_14076_ _03921_ _03942_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__nor2_1
X_11288_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[105\] _07111_
+ _07130_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[97\] vssd1 vssd1
+ vccd1 vccd1 _07248_ sky130_fd_sc_hd__a22o_1
X_17904_ clknet_leaf_90_wb_clk_i _03247_ _01600_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08338__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13027_ net305 net2763 net461 vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__mux2_1
X_10239_ _05911_ net511 net336 _06263_ vssd1 vssd1 vccd1 vccd1 _06264_ sky130_fd_sc_hd__o22a_1
XANTENNA_clkbuf_leaf_67_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10143__A _04490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1040 team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[23\]
+ vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09491__X team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1051 net1065 vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__buf_4
XFILLER_0_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17835_ clknet_leaf_74_wb_clk_i _03178_ _01531_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[81\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1062 net1063 vssd1 vssd1 vccd1 vccd1 net1062 sky130_fd_sc_hd__buf_4
XANTENNA__12769__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1073 net1076 vssd1 vssd1 vccd1 vccd1 net1073 sky130_fd_sc_hd__buf_4
XFILLER_0_156_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1084 net1086 vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__buf_4
XANTENNA__17571__D team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1095 net1097 vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__buf_4
XANTENNA__09651__B net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17766_ clknet_leaf_84_wb_clk_i _03109_ _01462_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_14978_ net1204 vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16717_ clknet_leaf_159_wb_clk_i _02347_ _00413_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13929_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[2\] team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[1\]
+ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[3\] vssd1 vssd1 vccd1
+ vccd1 _03804_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11645__A2 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17697_ clknet_leaf_98_wb_clk_i _03040_ _01393_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[71\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08510__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16648_ clknet_leaf_204_wb_clk_i _02278_ _00344_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14285__A _06424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16579_ clknet_leaf_198_wb_clk_i _02209_ _00275_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_09120_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[12\]
+ net837 net755 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_106_Left_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18318_ net1410 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_44_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09051_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[13\]
+ net672 net656 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__a22o_1
X_18249_ clknet_leaf_38_wb_clk_i _03478_ _01944_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_115_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09223__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold501 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1915 sky130_fd_sc_hd__dlygate4sd3_1
Xhold512 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[6\] vssd1
+ vssd1 vccd1 vccd1 net1926 sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 team_05_WB.instance_to_wrap.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 net1937
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08577__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold534 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 net1948 sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1959 sky130_fd_sc_hd__dlygate4sd3_1
Xhold556 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[68\] vssd1 vssd1
+ vccd1 vccd1 net1970 sky130_fd_sc_hd__dlygate4sd3_1
Xhold567 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net1981 sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net1992 sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ _05981_ vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__inv_2
Xhold589 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2003 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_115_Left_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08904_ _04944_ _04966_ vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__and2b_1
X_09884_ _04594_ _05912_ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout1107_A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1201 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net2615 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1212 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2626 sky130_fd_sc_hd__dlygate4sd3_1
X_08835_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[18\]
+ net810 _04406_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__a22o_1
Xhold1223 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2637 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1234 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2648 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11436__X _07349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout567_A _06774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1245 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net2659 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1256 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2670 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1267 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2681 sky130_fd_sc_hd__dlygate4sd3_1
X_08766_ _04824_ _04837_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[21\]
+ net592 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[21\]
+ sky130_fd_sc_hd__o2bb2a_4
Xhold1278 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 net2692 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09829__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1289 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2703 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11155__Y _07121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08697_ _04763_ _04765_ _04767_ _04769_ vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__or4_2
XFILLER_0_67_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout734_A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout901_A net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout522_X net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13303__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09318_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[8\]
+ net797 _05361_ vssd1 vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_157_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10590_ net1020 _05281_ _05283_ net551 vssd1 vssd1 vccd1 vccd1 _06598_ sky130_fd_sc_hd__a211o_1
XANTENNA__12061__A2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[12\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09249_ _05295_ _05297_ _05298_ _05299_ vssd1 vssd1 vccd1 vccd1 _05300_ sky130_fd_sc_hd__or4_1
XFILLER_0_17_972 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12260_ _07963_ _07964_ _07966_ _03554_ vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__a211o_1
XANTENNA__09214__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout891_X net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11211_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[109\] _07111_
+ _07125_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[21\] _07174_
+ vssd1 vssd1 vccd1 vccd1 _07175_ sky130_fd_sc_hd__a221o_1
XFILLER_0_105_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_101_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08568__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12191_ _08001_ _08002_ vssd1 vssd1 vccd1 vccd1 _08003_ sky130_fd_sc_hd__nand2_1
XANTENNA__11572__B2 _07396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11142_ _07072_ _07107_ vssd1 vssd1 vccd1 vccd1 _07108_ sky130_fd_sc_hd__nor2_4
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__clkbuf_4
XANTENNA__09517__A1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[10\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__clkbuf_4
X_11073_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[3\] _07035_
+ _04161_ _04162_ vssd1 vssd1 vccd1 vccd1 _07040_ sky130_fd_sc_hd__a211o_1
X_15950_ net1272 vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 ADR_O[30] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input30_A DAT_I[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14901_ net1060 vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__inv_2
X_10024_ net1020 _04427_ net553 _04426_ vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__a211o_1
XANTENNA__12589__S net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15881_ net1276 vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__inv_2
X_17620_ clknet_leaf_58_wb_clk_i _02991_ _01316_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08740__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14832_ net1183 vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_172_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_172_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17551_ clknet_leaf_57_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[22\]
+ _01247_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[22\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_101_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_101_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_14763_ net1070 vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__inv_2
X_11975_ _07749_ _07777_ _07785_ _07719_ vssd1 vssd1 vccd1 vccd1 _07787_ sky130_fd_sc_hd__a31o_1
XANTENNA_output117_A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16502_ clknet_leaf_142_wb_clk_i _02132_ _00198_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13714_ net899 _06521_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[14\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10926_ _05900_ _05905_ vssd1 vssd1 vccd1 vccd1 _06917_ sky130_fd_sc_hd__nor2_1
X_17482_ clknet_leaf_26_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[17\]
+ _01178_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14694_ net1208 vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__inv_2
X_16433_ clknet_leaf_118_wb_clk_i _02063_ _00129_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13721__B _06387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10857_ _06852_ _06853_ _06827_ vssd1 vssd1 vccd1 vccd1 _06854_ sky130_fd_sc_hd__a21bo_1
X_13645_ net2766 net278 net388 vssd1 vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__mux2_1
XANTENNA__12588__A0 _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13213__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_140_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16364_ clknet_leaf_2_wb_clk_i _01994_ _00060_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10788_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[26\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06785_ sky130_fd_sc_hd__or2_1
X_13576_ net2896 net271 net396 vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09453__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18103_ clknet_leaf_52_wb_clk_i _03426_ _01799_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11260__B1 _07124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15315_ net1214 vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14329__A1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12527_ _07812_ net1842 _03675_ vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16295_ net1143 vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18034_ clknet_leaf_97_wb_clk_i _03373_ _01730_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15246_ net1179 vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__inv_2
XFILLER_0_169_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12458_ net1689 _07812_ _03670_ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__mux2_1
XANTENNA__17917__Q team_05_WB.instance_to_wrap.wishbone.curr_state\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11409_ net2219 _07327_ vssd1 vssd1 vccd1 vccd1 _07335_ sky130_fd_sc_hd__nor2_1
X_12389_ net1673 _03664_ net216 vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__mux2_1
XANTENNA__10425__X _06442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15177_ net1221 vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__inv_2
XANTENNA__09646__B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14128_ _03803_ _03984_ _03987_ _03990_ _03858_ vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__a41o_1
XFILLER_0_123_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14059_ _03905_ _03907_ _03926_ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__nand3_1
XFILLER_0_94_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wire535_A _05234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12499__S net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08620_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[24\]
+ net684 net677 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[24\]
+ _04680_ vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__a221o_1
X_17818_ clknet_leaf_102_wb_clk_i _03161_ _01514_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[64\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08731__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08551_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[26\]
+ net804 net773 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__a22o_1
X_17749_ clknet_leaf_92_wb_clk_i _03092_ _01445_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08482_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[27\]
+ net696 net677 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[27\]
+ _04555_ vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_46_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12579__A0 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13123__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11432__A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12043__A2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[25\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09103_ _05153_ _05155_ _05157_ _05159_ vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_135_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11251__B1 _07121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08798__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10048__A _04656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout315_A net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09034_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[14\]
+ net803 net789 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11003__B1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold320 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[109\] vssd1 vssd1
+ vccd1 vccd1 net1734 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold331 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[127\] vssd1 vssd1
+ vccd1 vccd1 net1745 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold342 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[72\] vssd1 vssd1
+ vccd1 vccd1 net1756 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1224_A net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold353 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[90\] vssd1 vssd1
+ vccd1 vccd1 net1767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 net95 vssd1 vssd1 vccd1 vccd1 net1778 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold375 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[32\] vssd1 vssd1
+ vccd1 vccd1 net1789 sky130_fd_sc_hd__dlygate4sd3_1
Xhold386 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[44\] vssd1 vssd1
+ vccd1 vccd1 net1800 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout684_A net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout800 net801 vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__buf_4
Xhold397 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[112\] vssd1 vssd1
+ vccd1 vccd1 net1811 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout811 net813 vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_68_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09936_ _05104_ _05935_ vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__nor2_1
Xfanout822 net825 vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1012_X net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout833 net836 vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__clkbuf_8
Xfanout844 _04375_ vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__buf_4
Xfanout855 _04367_ vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__clkbuf_8
Xfanout866 _04291_ vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17562__Q team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09867_ net379 _04716_ vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout851_A _04370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout877 net882 vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__buf_1
XANTENNA_fanout472_X net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout888 _04280_ vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__clkbuf_4
Xhold1020 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net2434 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout899 _04235_ vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__clkbuf_4
Xhold1031 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2445 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout949_A _04363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1042 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2456 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08722__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1053 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2467 sky130_fd_sc_hd__dlygate4sd3_1
X_08818_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[18\]
+ net707 net656 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__a22o_1
XFILLER_0_169_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09798_ _05188_ _05828_ _05186_ vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__a21o_2
Xhold1064 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2478 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09722__D net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1075 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net2489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1086 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 net2500 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1097 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 net2511 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08749_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[21\]
+ net838 net779 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout737_X net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _07569_ _07571_ vssd1 vssd1 vccd1 vccd1 _07572_ sky130_fd_sc_hd__and2_1
XFILLER_0_166_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10293__A1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[25\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10711_ _06711_ _06710_ _06646_ net525 vssd1 vssd1 vccd1 vccd1 _06712_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10293__B2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[25\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11691_ net913 vssd1 vssd1 vccd1 vccd1 _07504_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout904_X net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13033__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13430_ net1950 net189 net413 vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__mux2_1
X_10642_ net529 _06646_ net335 vssd1 vssd1 vccd1 vccd1 _06647_ sky130_fd_sc_hd__a21o_1
XANTENNA__09435__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11242__B1 _07105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_5_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13361_ net557 _03694_ _03701_ vssd1 vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__and3_1
XANTENNA__12872__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10573_ _06505_ _06581_ net529 vssd1 vssd1 vccd1 vccd1 _06582_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_172_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15100_ net1097 vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12312_ _03604_ _03605_ _03606_ vssd1 vssd1 vccd1 vccd1 _03607_ sky130_fd_sc_hd__nand3_1
X_16080_ net1259 vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13292_ net322 net2649 net432 vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09738__A1 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12243_ net355 _03518_ vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15031_ net1097 vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__inv_2
XANTENNA__10245__X _06270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12742__A0 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12174_ _07982_ _07983_ _07985_ vssd1 vssd1 vccd1 vccd1 _07986_ sky130_fd_sc_hd__a21oi_2
XANTENNA__10405__B _06422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11125_ _07081_ _07087_ vssd1 vssd1 vccd1 vccd1 _07091_ sky130_fd_sc_hd__nor2_4
X_16982_ clknet_leaf_142_wb_clk_i _02612_ _00678_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11056_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[11\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[10\]
+ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[13\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[12\]
+ vssd1 vssd1 vccd1 vccd1 _07023_ sky130_fd_sc_hd__or4_1
X_15933_ net1269 vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__inv_2
XANTENNA__13716__B _06481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17472__Q team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[7\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08713__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13208__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10007_ _06034_ _06035_ vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__nand2_1
X_15864_ net1265 vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__inv_2
X_17603_ clknet_leaf_80_wb_clk_i _02974_ _01299_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_14815_ net1180 vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15795_ net1305 vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17534_ clknet_leaf_80_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[5\]
+ _01230_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13732__A net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14746_ net1052 vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__inv_2
X_11958_ _07767_ _07769_ vssd1 vssd1 vccd1 vccd1 _07770_ sky130_fd_sc_hd__nor2_1
XANTENNA__08385__X team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[30\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10909_ _06781_ _06783_ _06882_ net1044 vssd1 vssd1 vccd1 vccd1 _06903_ sky130_fd_sc_hd__o31a_1
X_17465_ clknet_leaf_36_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[0\]
+ _01161_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14677_ net1079 vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11889_ _07699_ _07700_ vssd1 vssd1 vccd1 vccd1 _07701_ sky130_fd_sc_hd__nor2_1
XANTENNA__11252__A _07031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16416_ clknet_leaf_131_wb_clk_i _02046_ _00112_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13628_ net2659 net190 net389 vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__mux2_1
X_17396_ clknet_leaf_60_wb_clk_i net1436 _01092_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09426__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13222__A1 _06687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11233__B1 _07119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16347_ clknet_leaf_191_wb_clk_i _01977_ _00043_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12782__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13559_ _04252_ net557 _03707_ vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__and3_4
XFILLER_0_82_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12981__A0 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16278_ net1158 vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14282__B _06591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18017_ clknet_leaf_82_wb_clk_i _03356_ _01713_ vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_130_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15229_ net1090 vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__inv_2
XANTENNA__10155__X _06183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08280__B team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[21\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12733__A0 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09721_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[0\]
+ net1017 net951 net926 vssd1 vssd1 vccd1 vccd1 _05753_ sky130_fd_sc_hd__and4_1
XANTENNA__10602__Y _06609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13118__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08704__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09652_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[1\]
+ net940 net932 net930 vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__and4_1
X_08603_ _04677_ vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__inv_2
X_09583_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[2\]
+ net940 net930 net927 vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__and4_1
XANTENNA__12957__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08534_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[26\]
+ net631 _04610_ net722 vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__a211o_1
XFILLER_0_89_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09665__B1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08465_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[28\]
+ net824 net797 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[28\]
+ _04543_ vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout432_A _03722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1174_A net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_154_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08396_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[29\]
+ net619 net599 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__a22o_1
XFILLER_0_163_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14473__A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_150_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10983__C1 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_947 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout899_A _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09017_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[14\]
+ net718 _05072_ _05077_ vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__o22a_4
XFILLER_0_14_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_783 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09717__D _04418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold150 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[9\]
+ vssd1 vssd1 vccd1 vccd1 net1564 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09196__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold161 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[14\]
+ vssd1 vssd1 vccd1 vccd1 net1575 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[31\]
+ vssd1 vssd1 vccd1 vccd1 net1586 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold183 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[21\]
+ vssd1 vssd1 vccd1 vccd1 net1597 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout687_X net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold194 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[27\] vssd1 vssd1
+ vccd1 vccd1 net1608 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08943__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout630 net631 vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__clkbuf_8
Xfanout641 net643 vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_109_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout652 net655 vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__buf_6
X_09919_ _05669_ _05946_ _05943_ vssd1 vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_109_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout663 _04306_ vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__buf_4
Xfanout674 net675 vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__buf_4
XANTENNA_fanout854_X net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout685 net686 vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__clkbuf_8
X_12930_ net197 net2435 net469 vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout696 net698 vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_126_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_126_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12867__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12861_ net562 _03698_ _03702_ vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__or3_1
XANTENNA__09105__C1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14600_ net1218 vssd1 vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__inv_2
X_11812_ _07602_ _07607_ _07609_ vssd1 vssd1 vccd1 vccd1 _07624_ sky130_fd_sc_hd__and3_1
X_15580_ net1250 vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12792_ net307 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[0\]
+ net489 vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09120__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14531_ net1196 vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__inv_2
X_11743_ _07545_ _07550_ _07546_ _07532_ vssd1 vssd1 vccd1 vccd1 _07555_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10387__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17250_ clknet_leaf_7_wb_clk_i _02880_ _00946_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09408__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14462_ net1062 vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11674_ _04167_ _07486_ net1049 net507 vssd1 vssd1 vccd1 vccd1 _07489_ sky130_fd_sc_hd__or4b_1
XFILLER_0_126_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16201_ net1110 vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__inv_2
XANTENNA__11215__B1 _07126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13413_ net2749 net282 net417 vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10625_ _05378_ _06056_ vssd1 vssd1 vccd1 vccd1 _06631_ sky130_fd_sc_hd__nand2_1
X_17181_ clknet_leaf_111_wb_clk_i _02811_ _00877_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_14393_ net1553 vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16132_ net1277 vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__inv_2
X_10556_ _06049_ _06229_ _06558_ net554 vssd1 vssd1 vccd1 vccd1 _06566_ sky130_fd_sc_hd__o22a_1
X_13344_ net268 net2393 net424 vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16063_ net1262 vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__inv_2
X_10487_ _05835_ _05935_ vssd1 vssd1 vccd1 vccd1 _06500_ sky130_fd_sc_hd__xnor2_4
X_13275_ net257 net2144 net433 vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__mux2_1
XANTENNA__11518__A1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11011__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09187__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15014_ net1247 vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__inv_2
X_12226_ _08016_ _08019_ _08017_ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08395__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13727__A net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12157_ _07963_ _07964_ _07966_ vssd1 vssd1 vccd1 vccd1 _07969_ sky130_fd_sc_hd__a21o_2
XANTENNA__08934__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16103__A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11108_ _07063_ _07067_ vssd1 vssd1 vccd1 vccd1 _07075_ sky130_fd_sc_hd__and2b_2
XFILLER_0_120_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16965_ clknet_leaf_19_wb_clk_i _02595_ _00661_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12088_ _07886_ _07887_ _07899_ _07888_ vssd1 vssd1 vccd1 vccd1 _07900_ sky130_fd_sc_hd__o31a_1
XANTENNA__09643__C net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15916_ net1305 vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__inv_2
X_11039_ _07009_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[5\] net569
+ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_34_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16896_ clknet_leaf_132_wb_clk_i _02526_ _00592_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_15847_ net1293 vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__inv_2
XANTENNA__12777__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14558__A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15778_ net1297 vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10257__A1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17517_ clknet_leaf_74_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[20\]
+ _01213_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09111__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14729_ net1222 vssd1 vssd1 vccd1 vccd1 _00359_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08250_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[31\]
+ net622 net615 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__a22o_1
X_17448_ clknet_leaf_50_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[16\]
+ _01144_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11206__B1 _07124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08181_ _04258_ _04263_ vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__and2_4
X_17379_ clknet_leaf_81_wb_clk_i net1437 _01075_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12365__X _03660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14293__A _04573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_9_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13401__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08291__A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13903__C1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09178__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_204_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_204_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_58_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_151_Right_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09851__A_N net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout382_A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09704_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[20\] _04267_
+ _05212_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[7\] _05736_
+ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[0\]
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_65_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11693__A0 team_05_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09635_ net954 _04267_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__o21a_1
XANTENNA__09350__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1291_A net1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09566_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[2\]
+ net1015 net947 net924 vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__and4_1
XANTENNA__09102__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08517_ _04573_ _04593_ vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__or2_1
X_09497_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[4\]
+ net618 net615 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[4\]
+ _05535_ vssd1 vssd1 vccd1 vccd1 _05536_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout814_A _04388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout435_X net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1177_X net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08310__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08448_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[28\]
+ net667 net662 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13198__A0 _06270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08379_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[30\]
+ net758 net739 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[30\]
+ _04459_ vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout602_X net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10410_ net888 _05974_ _06426_ vssd1 vssd1 vccd1 vccd1 _06427_ sky130_fd_sc_hd__or3_1
XANTENNA__13311__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwire349 _05305_ vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__buf_4
X_11390_ _07315_ net730 vssd1 vssd1 vccd1 vccd1 _07321_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10956__C1 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10341_ _06353_ _06356_ _06361_ net537 vssd1 vssd1 vccd1 vccd1 _06362_ sky130_fd_sc_hd__a31o_1
XANTENNA__09169__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13060_ net305 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[0\]
+ net456 vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__mux2_1
X_10272_ _05900_ _05989_ net894 vssd1 vssd1 vccd1 vccd1 _06295_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12011_ net343 _07691_ vssd1 vssd1 vccd1 vccd1 _07823_ sky130_fd_sc_hd__nor2_1
XANTENNA__08377__B1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08916__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout460 _03711_ vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__buf_6
Xfanout471 _03709_ vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__clkbuf_8
Xfanout482 net483 vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__buf_8
X_16750_ clknet_leaf_171_wb_clk_i _02380_ _00446_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13962_ _03816_ _03833_ vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_6_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout493 _03699_ vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__buf_4
XANTENNA__08928__X team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[16\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13673__A1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15701_ net1152 vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_79_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09341__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12913_ net284 net2753 net473 vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__mux2_1
XANTENNA__12597__S _03680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16681_ clknet_leaf_18_wb_clk_i _02311_ _00377_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13893_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[18\]
+ net558 net574 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[18\]
+ net985 vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__a221o_1
X_15632_ net1248 vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__inv_2
X_12844_ net267 net2966 net480 vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18351_ net1336 vssd1 vssd1 vccd1 vccd1 irq[2] sky130_fd_sc_hd__buf_2
XANTENNA__10239__B2 _06263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15563_ net1246 vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__inv_2
X_12775_ net261 net2734 net488 vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__mux2_1
X_17302_ clknet_leaf_151_wb_clk_i _02932_ _00998_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14514_ net1239 vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18282_ net107 vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__clkbuf_1
X_11726_ _07379_ _07447_ _07536_ vssd1 vssd1 vccd1 vccd1 _07538_ sky130_fd_sc_hd__or3_1
X_15494_ net1158 vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_778 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17233_ clknet_leaf_122_wb_clk_i _02863_ _00929_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14445_ net1081 vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__inv_2
X_11657_ net5 net990 net917 net1547 vssd1 vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__o22a_1
XFILLER_0_153_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10608_ net1020 _05331_ net553 vssd1 vssd1 vccd1 vccd1 _06615_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17164_ clknet_leaf_0_wb_clk_i _02794_ _00860_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_14376_ _04168_ net1542 _07451_ vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__a21o_1
X_11588_ _07354_ _07384_ net546 net1007 net75 vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__a32o_1
XANTENNA__09638__C net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16115_ net1134 vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold908 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2322 sky130_fd_sc_hd__dlygate4sd3_1
X_13327_ net2037 net306 net431 vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__mux2_1
X_10539_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[12\] _06091_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06550_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08080__A2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[21\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold919 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2333 sky130_fd_sc_hd__dlygate4sd3_1
X_17095_ clknet_leaf_200_wb_clk_i _02725_ _00791_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10146__A _04573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10962__A2 _06768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16046_ net1251 vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__inv_2
X_13258_ net309 net2289 net436 vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__mux2_1
XANTENNA__08368__B1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12209_ _08014_ _08018_ _08020_ _08012_ _08009_ vssd1 vssd1 vccd1 vccd1 _08021_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08907__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10580__S net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13900__A2 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13189_ net309 net2738 net441 vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__mux2_1
XANTENNA__11372__C1 _06769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17997_ clknet_leaf_83_wb_clk_i _03336_ _01693_ vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__dfrtp_1
XANTENNA__13113__A0 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16948_ clknet_leaf_115_wb_clk_i _02578_ _00644_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_84_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09332__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16879_ clknet_leaf_137_wb_clk_i _02509_ _00575_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14288__A _06219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08540__B1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09420_ net573 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[6\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[6\] vssd1 vssd1 vccd1
+ vccd1 _05463_ sky130_fd_sc_hd__a21oi_1
X_09351_ net953 _04350_ _04269_ vssd1 vssd1 vccd1 vccd1 _05398_ sky130_fd_sc_hd__a21o_1
XANTENNA__13967__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08302_ net1016 net943 net933 vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__and3_1
XFILLER_0_157_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09282_ net349 _05329_ vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08233_ net884 net865 net861 vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10755__S net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13131__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14335__A2_N net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08164_ net956 _04246_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__nand2_2
XFILLER_0_15_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08095_ net1027 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__and2b_1
XANTENNA__12970__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10056__A team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1137_A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload70 clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload70/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_113_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload81 clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload81/Y sky130_fd_sc_hd__inv_6
Xclkload92 clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload92/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__08359__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11439__X _07352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09020__A1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[26\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09564__B net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11158__Y _07124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout385_X net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout764_A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08997_ _05034_ _05055_ vssd1 vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09323__A2 _04366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout552_X net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08531__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13306__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09618_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[2\]
+ net880 net870 _04289_ vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__and4_1
X_10890_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[31\] net1041 vssd1
+ vssd1 vccd1 vccd1 _06887_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09087__A1 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09549_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[3\]
+ net712 net598 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[3\]
+ _05578_ vssd1 vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout817_X net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12560_ _03632_ net1847 net207 vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08834__A1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[30\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11511_ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[20\] _07421_ net1003
+ vssd1 vssd1 vccd1 vccd1 _07422_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_197_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_197_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12491_ net1626 _03632_ net210 vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__mux2_1
XANTENNA__09897__A_N net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13041__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14230_ team_05_WB.instance_to_wrap.total_design.keypad0.counter\[15\] _04025_ vssd1
+ vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11442_ net920 _07354_ vssd1 vssd1 vccd1 vccd1 _07355_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_126_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_126_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11197__A2 _07128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11373_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[0\] _06769_ _07310_
+ vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__o21ba_1
X_14161_ _03970_ net907 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[10\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__12880__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08062__A2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[30\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input60_A wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10324_ _06342_ _06345_ _04265_ vssd1 vssd1 vccd1 vccd1 _06346_ sky130_fd_sc_hd__o21a_2
X_13112_ net277 net2641 net450 vssd1 vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__mux2_1
X_14092_ _03940_ _03957_ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11496__S net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13343__A0 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17920_ clknet_leaf_35_wb_clk_i _03259_ _01616_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10255_ _06277_ _06278_ net370 vssd1 vssd1 vccd1 vccd1 _06279_ sky130_fd_sc_hd__mux2_1
X_13043_ net259 net2696 net457 vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_57_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_147_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1200 net1202 vssd1 vssd1 vccd1 vccd1 net1200 sky130_fd_sc_hd__buf_4
Xfanout1211 net1313 vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__clkbuf_4
X_17851_ clknet_leaf_75_wb_clk_i _03194_ _01547_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[33\]
+ sky130_fd_sc_hd__dfrtp_1
X_10186_ _06189_ _06204_ _06212_ net537 vssd1 vssd1 vccd1 vccd1 _06213_ sky130_fd_sc_hd__a31o_1
Xfanout1222 net1225 vssd1 vssd1 vccd1 vccd1 net1222 sky130_fd_sc_hd__buf_4
Xfanout1233 net1234 vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__buf_4
Xfanout1244 net1252 vssd1 vssd1 vccd1 vccd1 net1244 sky130_fd_sc_hd__buf_4
Xfanout1255 net1279 vssd1 vssd1 vccd1 vccd1 net1255 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08770__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16802_ clknet_leaf_15_wb_clk_i _02432_ _00498_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_17782_ clknet_leaf_88_wb_clk_i _03125_ _01478_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[28\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1266 net1268 vssd1 vssd1 vccd1 vccd1 net1266 sky130_fd_sc_hd__buf_2
Xfanout1277 net1278 vssd1 vssd1 vccd1 vccd1 net1277 sky130_fd_sc_hd__buf_2
X_14994_ net1235 vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1288 net1291 vssd1 vssd1 vccd1 vccd1 net1288 sky130_fd_sc_hd__buf_4
Xfanout290 net293 vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__clkbuf_2
Xfanout1299 net1300 vssd1 vssd1 vccd1 vccd1 net1299 sky130_fd_sc_hd__buf_4
XANTENNA__09314__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16733_ clknet_leaf_108_wb_clk_i _02363_ _00429_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13724__B _06320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13945_ _03810_ _03818_ _07451_ vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__o21a_1
XFILLER_0_89_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13216__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08522__B1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload6_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16664_ clknet_leaf_30_wb_clk_i _02294_ _00360_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13876_ net1564 net983 _03774_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[9\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_72_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09640__D net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15615_ net1156 vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__inv_2
X_18403_ net1373 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__buf_2
X_12827_ net308 net2855 net484 vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__mux2_1
X_16595_ clknet_leaf_154_wb_clk_i _02225_ _00291_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18334_ net1323 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
XFILLER_0_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15546_ net1123 vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12758_ net324 net2944 net493 vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17569__D team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18265_ clknet_leaf_36_wb_clk_i _03494_ _01960_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[19\]
+ sky130_fd_sc_hd__dfrtp_4
X_11709_ _07476_ _07520_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[4\]
+ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[5\] vssd1 vssd1 vccd1
+ vccd1 _07521_ sky130_fd_sc_hd__or4bb_1
X_15477_ net1172 vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12689_ net1976 net340 vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__and2_1
XFILLER_0_142_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17216_ clknet_leaf_132_wb_clk_i _02846_ _00912_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14428_ net1074 vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18196_ clknet_leaf_37_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[17\]
+ _01891_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11188__A2 _07105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12385__A1 _07812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08589__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_96_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_170_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17147_ clknet_leaf_191_wb_clk_i _02777_ _00843_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold705 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 net2119 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12790__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14359_ _04109_ _04108_ vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__nand2b_1
XANTENNA__10396__B1 _06055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold716 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net2141 sky130_fd_sc_hd__dlygate4sd3_1
Xhold738 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2152 sky130_fd_sc_hd__dlygate4sd3_1
X_17078_ clknet_leaf_150_wb_clk_i _02708_ _00774_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold749 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net2163 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08920_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[16\]
+ net621 net602 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16029_ net1285 vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09553__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08851_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[18\]
+ net778 net764 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[18\]
+ _04905_ vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_51_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1405 _03291_ vssd1 vssd1 vccd1 vccd1 net2819 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08761__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1416 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2830 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1427 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 net2841 sky130_fd_sc_hd__dlygate4sd3_1
X_08782_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[19\]
+ net711 net698 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[19\]
+ _04852_ vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__a221o_1
Xhold1438 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 net2852 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1449 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2863 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13193__Y _03717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_203_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13126__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09403_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[6\]
+ net833 net794 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_49_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12965__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout345_A net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1087_A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09334_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[7\]
+ net645 net600 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[7\]
+ _05379_ vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11441__Y _07354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09265_ _05313_ _05314_ vssd1 vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout512_A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08216_ net879 net862 net858 vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09196_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[10\]
+ net644 net598 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[10\]
+ _05248_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12376__A1 _03646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11179__A2 _07092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08147_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[3\] team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[2\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[1\] team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__and4bb_2
XTAP_TAPCELL_ROW_116_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload170 clknet_leaf_88_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload170/Y sky130_fd_sc_hd__bufinv_16
X_08078_ net1023 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[22\]
+ net970 _04188_ vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__a22o_1
Xclkload181 clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload181/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_141_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout881_A net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload192 clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload192/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_112_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10514__A _06525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10040_ _06067_ _06068_ vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_164_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09544__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold10 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[13\]
+ vssd1 vssd1 vccd1 vccd1 net1424 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[25\]
+ vssd1 vssd1 vccd1 vccd1 net1435 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout767_X net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold32 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1446 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[16\] vssd1 vssd1
+ vccd1 vccd1 net1457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[5\]
+ vssd1 vssd1 vccd1 vccd1 net1468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[24\] vssd1 vssd1
+ vccd1 vccd1 net1479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[22\]
+ vssd1 vssd1 vccd1 vccd1 net1490 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[29\]
+ vssd1 vssd1 vccd1 vccd1 net1501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[26\] vssd1 vssd1
+ vccd1 vccd1 net1512 sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ net356 _07538_ _07784_ _07796_ vssd1 vssd1 vccd1 vccd1 _07803_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_97_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout934_X net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09741__C net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08197__Y _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08504__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13036__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13730_ net899 _06108_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[30\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10942_ _06927_ _06930_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[23\]
+ net564 vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_168_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13661_ net2017 net190 net386 vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__mux2_1
X_10873_ _06802_ _06869_ vssd1 vssd1 vccd1 vccd1 _06870_ sky130_fd_sc_hd__nand2_1
XANTENNA__12875__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15400_ net1224 vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__inv_2
X_12612_ _07367_ _07859_ _07863_ _03659_ vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__or4b_4
X_16380_ clknet_leaf_154_wb_clk_i _02010_ _00076_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_130_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13592_ _04250_ _04251_ _04256_ net557 vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__and4_4
XFILLER_0_38_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15331_ net1197 vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__inv_2
X_12543_ _07840_ _07851_ _03677_ vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__and3_4
XFILLER_0_136_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18050_ net1039 _03388_ _01746_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_124_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15262_ net1066 vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__inv_2
X_12474_ _07840_ _07850_ _03672_ vssd1 vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__and3_4
XFILLER_0_35_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12367__A1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[30\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10408__B _06424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17001_ clknet_leaf_15_wb_clk_i _02631_ _00697_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14213_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[12\] _04011_
+ vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13559__X _03731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11425_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[1\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[0\]
+ net2110 vssd1 vssd1 vccd1 vccd1 _07341_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15193_ net1053 vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__inv_2
XANTENNA_7 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14144_ net1624 net502 net911 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[27\]
+ sky130_fd_sc_hd__and3_1
X_11356_ _07286_ _07288_ _07292_ vssd1 vssd1 vccd1 vccd1 _07298_ sky130_fd_sc_hd__and3_1
XANTENNA__13719__B _06424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10307_ _06328_ vssd1 vssd1 vccd1 vccd1 _06329_ sky130_fd_sc_hd__inv_2
X_14075_ _03921_ _03942_ vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__and2_1
X_11287_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[113\] _07104_
+ _07125_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[17\] vssd1 vssd1
+ vccd1 vccd1 _07247_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_94_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_17903_ clknet_leaf_88_wb_clk_i _03246_ _01599_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09535__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13026_ net326 net2043 net461 vssd1 vssd1 vccd1 vccd1 _02615_ sky130_fd_sc_hd__mux2_1
X_10238_ _06262_ vssd1 vssd1 vccd1 vccd1 _06263_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_4_0__f_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09912__A_N net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1030 net1036 vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10143__B net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13735__A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1041 team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[23\]
+ vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_23_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_17834_ clknet_leaf_98_wb_clk_i _03177_ _01530_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[80\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1052 net1053 vssd1 vssd1 vccd1 vccd1 net1052 sky130_fd_sc_hd__buf_2
X_10169_ net521 _06058_ vssd1 vssd1 vccd1 vccd1 _06196_ sky130_fd_sc_hd__nor2_1
Xfanout1063 net1064 vssd1 vssd1 vccd1 vccd1 net1063 sky130_fd_sc_hd__buf_4
Xfanout1074 net1075 vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__buf_4
Xfanout1085 net1086 vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__buf_2
Xfanout1096 net1097 vssd1 vssd1 vccd1 vccd1 net1096 sky130_fd_sc_hd__buf_4
X_17765_ clknet_leaf_100_wb_clk_i _03108_ _01461_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_14977_ net1223 vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__inv_2
XANTENNA__09651__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13928_ net978 team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[13\] team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[15\]
+ vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_16_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16716_ clknet_leaf_0_wb_clk_i _02346_ _00412_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_17696_ clknet_leaf_93_wb_clk_i _03039_ _01392_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[70\]
+ sky130_fd_sc_hd__dfrtp_1
X_16647_ clknet_leaf_201_wb_clk_i _02277_ _00343_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13859_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[1\]
+ net560 net576 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[1\]
+ net987 vssd1 vssd1 vccd1 vccd1 _03766_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12785__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14566__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16578_ clknet_leaf_6_wb_clk_i _02208_ _00274_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14285__B _06445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15529_ net1157 vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18317_ net1409 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_79_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09050_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[13\]
+ net651 net605 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[13\]
+ _05108_ vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__a221o_1
X_18248_ clknet_leaf_38_wb_clk_i _03477_ _01943_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18179_ clknet_leaf_42_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[0\]
+ _01874_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold502 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[116\] vssd1 vssd1
+ vccd1 vccd1 net1916 sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[87\] vssd1 vssd1
+ vccd1 vccd1 net1927 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10908__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold524 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[62\] vssd1 vssd1
+ vccd1 vccd1 net1938 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold535 net78 vssd1 vssd1 vccd1 vccd1 net1949 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold546 net139 vssd1 vssd1 vccd1 vccd1 net1960 sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 net1971 sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net1982 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08982__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09952_ _04798_ _04799_ vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__and2b_1
Xhold579 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net1993 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10334__A _05577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08903_ _04967_ vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__inv_2
XANTENNA__09526__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09883_ _04634_ _05907_ _05911_ vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__o21bai_2
XANTENNA__12530__A1 _03604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08734__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1202 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2616 sky130_fd_sc_hd__dlygate4sd3_1
X_08834_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[30\] net965
+ net953 _04902_ _04345_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[18\]
+ sky130_fd_sc_hd__a221o_1
Xhold1213 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 net2627 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1002_A _07345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10649__A1_N team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1224 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1235 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net2649 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1246 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2660 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1257 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2671 sky130_fd_sc_hd__dlygate4sd3_1
X_08765_ _04826_ _04830_ _04836_ vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__nor3_1
XANTENNA_fanout462_A _03711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1268 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 net2682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1279 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2693 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14179__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08696_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[22\]
+ net627 net608 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[22\]
+ _04768_ vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_68_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12695__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14476__A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout348_X net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08474__A _04552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12597__A1 _03663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09317_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[8\]
+ net804 net780 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[8\]
+ _05357_ vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_118_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout515_X net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12061__A3 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09857__X _05886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09248_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[9\]
+ net662 net626 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__a22o_1
XANTENNA__14338__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12349__A1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[20\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09179_ _05229_ _05230_ _05231_ _05232_ vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__or4_2
XFILLER_0_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11210_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[109\] _07102_
+ _07130_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[101\] vssd1
+ vssd1 vccd1 vccd1 _07174_ sky130_fd_sc_hd__a22o_1
X_12190_ _07941_ _07986_ _07981_ vssd1 vssd1 vccd1 vccd1 _08002_ sky130_fd_sc_hd__or3b_1
XANTENNA__09765__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11141_ _07068_ _07093_ vssd1 vssd1 vccd1 vccd1 _07107_ sky130_fd_sc_hd__nand2_2
XANTENNA__18411__A net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__clkbuf_4
X_11072_ _07036_ _07037_ vssd1 vssd1 vccd1 vccd1 _07039_ sky130_fd_sc_hd__nand2_8
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__clkbuf_4
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 ADR_O[31] sky130_fd_sc_hd__clkbuf_4
XANTENNA__12521__A1 _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10023_ _04157_ _05923_ vssd1 vssd1 vccd1 vccd1 _06052_ sky130_fd_sc_hd__or2_1
X_14900_ net1067 vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__inv_2
X_15880_ net1265 vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__inv_2
X_14831_ net1286 vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input23_A DAT_I[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17550_ clknet_leaf_59_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[21\]
+ _01246_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14762_ net1116 vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__inv_2
X_11974_ _07766_ _07780_ _07782_ _07784_ vssd1 vssd1 vccd1 vccd1 _07786_ sky130_fd_sc_hd__nand4_1
XANTENNA__09150__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16501_ clknet_leaf_71_wb_clk_i _02131_ _00197_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13713_ net900 _06540_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[13\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10925_ _06916_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[26\] net565
+ vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__mux2_1
X_17481_ clknet_leaf_37_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[16\]
+ _01177_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_14693_ net1193 vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16432_ clknet_leaf_166_wb_clk_i _02062_ _00128_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_141_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_141_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13644_ net2604 net282 net388 vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10856_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[8\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[8\]
+ vssd1 vssd1 vccd1 vccd1 _06853_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16363_ clknet_leaf_185_wb_clk_i _01993_ _00059_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13575_ net2547 net269 net396 vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__mux2_1
XANTENNA__08256__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10787_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[26\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06784_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18102_ clknet_leaf_52_wb_clk_i _03425_ _01798_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15314_ net1239 vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__inv_2
X_12526_ net1711 _03645_ net208 vssd1 vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14329__A2 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16294_ net1148 vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18033_ clknet_leaf_97_wb_clk_i _03372_ _01729_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_978 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15245_ net1082 vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12457_ net1636 _03645_ _03671_ vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11408_ net1939 _07328_ vssd1 vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_10_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09756__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15176_ net1224 vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__inv_2
X_12388_ _07478_ _03616_ vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__or2_4
XANTENNA__09646__C net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12353__B _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08964__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14127_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[15\] team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[12\]
+ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_91_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11339_ _04215_ team_05_WB.instance_to_wrap.total_design.keypad0.next_rows\[0\] _04228_
+ vssd1 vssd1 vccd1 vccd1 _07294_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_1_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09508__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14058_ _03905_ _03907_ _03926_ vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__a21o_1
XANTENNA__17582__D team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[19\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12512__A1 _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11315__A2 _07123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08716__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13009_ net263 net2256 net460 vssd1 vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__mux2_1
XANTENNA__08559__A _04613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08192__A1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17817_ clknet_leaf_100_wb_clk_i _03160_ _01513_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[127\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08550_ _04620_ _04622_ _04624_ _04626_ vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__or4_1
X_17748_ clknet_leaf_87_wb_clk_i _03091_ _01444_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09141__B1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08481_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[27\]
+ net680 net649 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[27\]
+ _04558_ vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_46_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17679_ clknet_leaf_88_wb_clk_i _03022_ _01375_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[117\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08495__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11713__A team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13404__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11432__B net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1056 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08247__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09102_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[12\]
+ net712 net695 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[12\]
+ _05158_ vssd1 vssd1 vccd1 vccd1 _05159_ sky130_fd_sc_hd__a221o_1
XANTENNA__10054__A2 _06033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09033_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[14\]
+ net811 net753 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[14\]
+ _05092_ vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__a221o_1
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout210_A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11003__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold310 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[87\] vssd1 vssd1
+ vccd1 vccd1 net1724 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold321 net130 vssd1 vssd1 vccd1 vccd1 net1735 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[70\] vssd1 vssd1
+ vccd1 vccd1 net1746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold343 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[91\] vssd1 vssd1
+ vccd1 vccd1 net1757 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08955__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold354 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[122\] vssd1 vssd1
+ vccd1 vccd1 net1768 sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[10\] vssd1 vssd1
+ vccd1 vccd1 net1779 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold376 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[61\] vssd1 vssd1
+ vccd1 vccd1 net1790 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold387 team_05_WB.instance_to_wrap.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1 net1801
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[26\]
+ vssd1 vssd1 vccd1 vccd1 net1812 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09853__A net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout801 _04394_ vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__buf_4
X_09935_ _05104_ _05963_ _05936_ vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__o21ai_1
Xfanout812 net813 vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__clkbuf_4
Xfanout823 net825 vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__clkbuf_8
Xfanout834 net836 vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12503__A1 _07816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11306__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout677_A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08707__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout845 _04373_ vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09572__B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout856 _04367_ vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__buf_4
X_09866_ net379 _04716_ vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__nor2_1
Xfanout867 net868 vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__buf_2
XANTENNA__13806__C net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1010 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2424 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout878 net879 vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__clkbuf_2
Xhold1021 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2435 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout889 _04280_ vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09380__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08817_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[18\]
+ net687 net602 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__a22o_1
Xhold1032 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2446 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1043 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 net2457 sky130_fd_sc_hd__dlygate4sd3_1
X_09797_ _05822_ _05827_ _05237_ vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__a21o_1
Xhold1054 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2468 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout844_A _04375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1065 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 net2479 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout465_X net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1076 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net2490 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08748_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[21\]
+ net799 net783 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__a22o_1
Xhold1087 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2501 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1098 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 net2512 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_2_0_wb_clk_i_X clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08486__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08679_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[23\]
+ net824 net739 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[23\]
+ _04740_ vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout632_X net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13314__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10710_ net517 _06006_ _06014_ net525 vssd1 vssd1 vccd1 vccd1 _06711_ sky130_fd_sc_hd__a31o_1
XANTENNA__10293__A2 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11690_ _07498_ _07499_ _07500_ _07503_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__or4_4
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10641_ _06611_ _06645_ net516 vssd1 vssd1 vccd1 vccd1 _06646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18406__A net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13360_ net306 net2072 net425 vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__mux2_1
X_10572_ _06543_ _06580_ net519 vssd1 vssd1 vccd1 vccd1 _06581_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_165_Right_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12311_ _07866_ _08022_ _03547_ _03603_ vssd1 vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__o22a_1
XFILLER_0_106_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13291_ net311 net2374 net433 vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15030_ net1091 vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__inv_2
X_12242_ _03524_ _03527_ _03512_ vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09738__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12173_ _07973_ _07975_ _07984_ _07977_ vssd1 vssd1 vccd1 vccd1 _07985_ sky130_fd_sc_hd__o31a_1
XFILLER_0_43_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08410__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11124_ net150 net732 vssd1 vssd1 vccd1 vccd1 _07090_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16981_ clknet_leaf_23_wb_clk_i _02611_ _00677_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15932_ net1305 vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__inv_2
X_11055_ _07022_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[2\] net566
+ vssd1 vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__mux2_1
XANTENNA__10505__B1 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09371__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10006_ net376 net364 vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__nand2_1
X_15863_ net1292 vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__inv_2
X_17602_ clknet_leaf_80_wb_clk_i _02973_ _01298_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_14814_ net1073 vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__inv_2
X_15794_ net1297 vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__inv_2
XANTENNA__09123__B1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17533_ clknet_leaf_81_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[4\]
+ _01229_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13732__B _06756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14745_ net1051 vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__inv_2
X_11957_ _07527_ _07752_ _07761_ vssd1 vssd1 vccd1 vccd1 _07769_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_28_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08477__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13224__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17464_ clknet_leaf_49_wb_clk_i net1050 _01160_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.last_read
+ sky130_fd_sc_hd__dfrtp_1
X_10908_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[29\] net568 _06902_
+ vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__a21o_1
X_14676_ net1074 vssd1 vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11888_ _07664_ _07669_ _07671_ vssd1 vssd1 vccd1 vccd1 _07700_ sky130_fd_sc_hd__and3_1
XFILLER_0_156_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16415_ clknet_leaf_156_wb_clk_i _02045_ _00111_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13627_ net2542 net195 net390 vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__mux2_1
X_17395_ clknet_leaf_65_wb_clk_i net1420 _01091_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_144_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10839_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[3\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06836_ sky130_fd_sc_hd__or2_1
XANTENNA__13222__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16346_ clknet_leaf_31_wb_clk_i _01976_ _00042_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13558_ net1945 net308 net401 vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_132_Right_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17577__D team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[14\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12509_ _07861_ _03659_ vssd1 vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__and2b_4
X_16277_ net1155 vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__inv_2
X_13489_ net312 net2324 net409 vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire380_A _04447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18016_ clknet_leaf_64_wb_clk_i _03355_ _01712_ vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__dfrtp_1
X_15228_ net1086 vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__inv_2
XANTENNA__09729__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08937__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15159_ net1102 vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__inv_2
XANTENNA__08401__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09720_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[0\]
+ net944 net939 net936 vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__and4_1
XANTENNA__09362__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09651_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[1\]
+ net1015 net946 net924 vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__and4_1
XFILLER_0_59_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08602_ _04656_ _04676_ vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__or2_1
XANTENNA__13923__A team_05_WB.instance_to_wrap.total_design.data_from_keypad\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09582_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[2\]
+ net947 net1013 net924 vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__and4_1
XANTENNA__09114__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08533_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[26\]
+ net681 net646 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08468__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout258_A _06442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13134__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_7_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08464_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[28\]
+ net835 net750 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_154_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12973__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08395_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[29\]
+ net711 net654 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__a22o_1
XFILLER_0_169_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout425_A _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1167_A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12421__A0 _03632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18309__1401 vssd1 vssd1 vccd1 vccd1 net1401 _18309__1401/LO sky130_fd_sc_hd__conb_1
XFILLER_0_18_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout213_X net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09016_ _05061_ _05074_ _05075_ _05076_ vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__or4_1
XFILLER_0_104_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout794_A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold140 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[17\] vssd1
+ vssd1 vccd1 vccd1 net1554 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[9\] vssd1 vssd1
+ vccd1 vccd1 net1565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[15\]
+ vssd1 vssd1 vccd1 vccd1 net1576 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10735__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold173 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[28\]
+ vssd1 vssd1 vccd1 vccd1 net1587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[18\]
+ vssd1 vssd1 vccd1 vccd1 net1598 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold195 team_05_WB.instance_to_wrap.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 net1609
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout961_A net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout582_X net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout620 _04317_ vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__buf_4
XANTENNA__13309__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout631 _04314_ vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__buf_6
Xfanout642 net643 vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__clkbuf_4
X_09918_ _05669_ _05946_ vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_109_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout653 net655 vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_109_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout664 _04305_ vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__buf_4
Xfanout675 _04303_ vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__buf_4
Xfanout686 _04300_ vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__buf_4
X_09849_ _04147_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[19\]
+ _04346_ _04359_ team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[21\]
+ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[20\]
+ sky130_fd_sc_hd__o41a_1
Xfanout697 net698 vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout847_X net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ net305 net2937 net480 vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__mux2_1
X_11811_ net549 _07622_ vssd1 vssd1 vccd1 vccd1 _07623_ sky130_fd_sc_hd__nand2_2
XFILLER_0_68_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10668__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12791_ net327 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[1\]
+ net489 vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__mux2_1
XANTENNA__08459__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13044__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ net1219 vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__inv_2
X_11742_ _07542_ _07547_ _07550_ _07553_ vssd1 vssd1 vccd1 vccd1 _07554_ sky130_fd_sc_hd__a211o_1
XFILLER_0_138_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14461_ net1090 vssd1 vssd1 vccd1 vccd1 _00091_ sky130_fd_sc_hd__inv_2
X_11673_ _07487_ vssd1 vssd1 vccd1 vccd1 _07488_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12883__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14664__A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16200_ net1146 vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12412__A0 _03657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13412_ net2031 net275 net419 vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17180_ clknet_leaf_158_wb_clk_i _02810_ _00876_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10624_ _06491_ net332 _06629_ net335 vssd1 vssd1 vccd1 vccd1 _06630_ sky130_fd_sc_hd__o22a_1
X_14392_ net1499 vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_133_Left_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16131_ net1277 vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13343_ net259 net2454 net425 vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10555_ net369 _06237_ net347 _06563_ _06564_ vssd1 vssd1 vccd1 vccd1 _06565_ sky130_fd_sc_hd__o311a_1
XANTENNA__10256__X _06280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08631__A2 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16062_ net1262 vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__inv_2
X_13274_ net254 net2500 net432 vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__mux2_1
X_10486_ net2085 net269 net539 vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11518__A2 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15013_ net1203 vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__inv_2
X_12225_ _03518_ _03519_ vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__nand2_1
XANTENNA__13727__B _06907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12156_ _07967_ _07963_ _07964_ vssd1 vssd1 vccd1 vccd1 _07968_ sky130_fd_sc_hd__mux2_2
XFILLER_0_166_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10703__Y _06705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11107_ _07073_ vssd1 vssd1 vccd1 vccd1 _07074_ sky130_fd_sc_hd__inv_2
XANTENNA__13219__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12087_ _07890_ _07885_ vssd1 vssd1 vccd1 vccd1 _07899_ sky130_fd_sc_hd__and2b_1
X_16964_ clknet_leaf_184_wb_clk_i _02594_ _00660_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09643__D _04418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_142_Left_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09344__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11038_ net964 _06672_ _07008_ vssd1 vssd1 vccd1 vccd1 _07009_ sky130_fd_sc_hd__a21oi_1
X_15915_ net1301 vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16895_ clknet_leaf_152_wb_clk_i _02525_ _00591_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08698__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13743__A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15846_ net1273 vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15777_ net1276 vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12989_ net314 net2901 net467 vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17516_ clknet_leaf_73_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[19\]
+ _01212_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_82_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12651__B1 _07349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14728_ net1218 vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17447_ clknet_leaf_60_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[15\]
+ _01143_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14659_ net1208 vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__inv_2
XANTENNA__14574__A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08870__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_151_Left_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08180_ _04261_ _04262_ vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__nor2_2
XFILLER_0_171_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17378_ clknet_leaf_81_wb_clk_i net1428 _01074_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14293__B team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[27\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09020__X team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[14\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16329_ net1125 vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__inv_2
XANTENNA__08622__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08291__B net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13903__B1 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08386__A1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_160_Left_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11438__A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13129__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09703_ net1019 net967 vssd1 vssd1 vccd1 vccd1 _05736_ sky130_fd_sc_hd__and2_1
XANTENNA__09335__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08689__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12968__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09634_ _05667_ _05668_ vssd1 vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__nand2_4
XFILLER_0_97_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09565_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[2\]
+ net947 net930 net925 vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout542_A _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08516_ _04592_ vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09496_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[4\]
+ net626 net608 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05535_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08447_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[28\]
+ net681 net596 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[28\]
+ _04525_ vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__a221o_1
XFILLER_0_147_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout428_X net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08861__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout807_A net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1072_X net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08378_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[30\]
+ net803 net742 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08613__A2 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10340_ _05924_ _06352_ _06360_ net348 vssd1 vssd1 vccd1 vccd1 _06361_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout797_X net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10271_ net2314 net242 net541 vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18289__1381 vssd1 vssd1 vccd1 vccd1 net1381 _18289__1381/LO sky130_fd_sc_hd__conb_1
XFILLER_0_104_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12010_ _07767_ _07769_ _07773_ _07774_ net549 vssd1 vssd1 vccd1 vccd1 _07822_ sky130_fd_sc_hd__o311a_1
XFILLER_0_104_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_47_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_40_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10523__Y _06535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout964_X net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09744__C net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13039__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout450 _03714_ vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__buf_6
Xfanout461 _03711_ vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__buf_4
Xfanout472 _03706_ vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__buf_6
X_13961_ _03816_ _03833_ vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__nor2_1
XANTENNA__12878__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout483 _03704_ vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__buf_4
Xfanout494 _03699_ vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__buf_6
X_15700_ net1152 vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__inv_2
X_12912_ net277 net2748 net475 vssd1 vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__mux2_1
X_16680_ clknet_leaf_203_wb_clk_i _02310_ _00376_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13892_ net1561 net981 _03782_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[17\]
+ sky130_fd_sc_hd__o21a_1
X_12843_ net260 net2399 net483 vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__mux2_1
X_15631_ net1246 vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18350_ net1335 vssd1 vssd1 vccd1 vccd1 irq[1] sky130_fd_sc_hd__buf_2
XANTENNA__12633__A0 _03604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15562_ net1131 vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__inv_2
XANTENNA__10239__A2 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12774_ net263 net2368 net488 vssd1 vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14513_ net1189 vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__inv_2
X_17301_ clknet_leaf_174_wb_clk_i _02931_ _00997_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_48_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11725_ _07379_ _07447_ _07478_ _07535_ vssd1 vssd1 vccd1 vccd1 _07537_ sky130_fd_sc_hd__or4_1
X_18281_ net107 vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__clkbuf_1
X_15493_ net1170 vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11811__A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13502__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17232_ clknet_leaf_152_wb_clk_i _02862_ _00928_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14444_ net1111 vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__inv_2
X_11656_ net6 net990 net917 net1577 vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__o22a_1
XFILLER_0_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17478__Q team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17163_ clknet_leaf_187_wb_clk_i _02793_ _00859_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10607_ _06469_ net332 _06613_ net335 vssd1 vssd1 vccd1 vccd1 _06614_ sky130_fd_sc_hd__o22a_1
XANTENNA_clkbuf_leaf_86_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14375_ net1039 _04043_ _00040_ vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11587_ _07354_ _07388_ net546 net1007 net1722 vssd1 vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__a32o_1
XANTENNA__08604__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16114_ net1135 vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__inv_2
XANTENNA__09638__D net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13326_ net1959 net324 net431 vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__mux2_1
Xhold909 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[17\] vssd1 vssd1
+ vccd1 vccd1 net2323 sky130_fd_sc_hd__dlygate4sd3_1
X_10538_ _06541_ _06542_ _06548_ _04275_ vssd1 vssd1 vccd1 vccd1 _06549_ sky130_fd_sc_hd__o31a_1
XFILLER_0_51_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17094_ clknet_leaf_115_wb_clk_i _02724_ _00790_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16045_ net1287 vssd1 vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__inv_2
XANTENNA__13738__A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13257_ net330 net2163 net438 vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10469_ net888 _05969_ _06482_ vssd1 vssd1 vccd1 vccd1 _06483_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12208_ _07999_ _08004_ _08006_ vssd1 vssd1 vccd1 vccd1 _08020_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_36_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13188_ net330 net2129 net442 vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12139_ _07943_ _07946_ _07948_ vssd1 vssd1 vccd1 vccd1 _07951_ sky130_fd_sc_hd__a21bo_1
X_17996_ clknet_leaf_83_wb_clk_i _03335_ _01692_ vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09317__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09951__A _05977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12788__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18308__1400 vssd1 vssd1 vccd1 vccd1 net1400 _18308__1400/LO sky130_fd_sc_hd__conb_1
X_16947_ clknet_leaf_168_wb_clk_i _02577_ _00643_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17590__D team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[27\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14569__A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09670__B net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16878_ clknet_leaf_177_wb_clk_i _02508_ _00574_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14288__B _06273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10910__A1_N net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15829_ net1256 vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08286__B _04366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12624__A0 _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09350_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[7\]
+ net717 _05392_ _05396_ vssd1 vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__o22ai_4
XANTENNA__09096__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08301_ net948 net1013 net927 vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__and3_2
XFILLER_0_75_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09281_ _05329_ vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08843__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13412__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09398__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[26\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08232_ net884 net875 net872 vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08163_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[3\] team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[1\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[0\] _04242_ vssd1
+ vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__nand4_4
XFILLER_0_67_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08094_ net1023 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[14\]
+ net970 _04196_ vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__a22o_1
XANTENNA__10056__B team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload60 clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload60/Y sky130_fd_sc_hd__inv_16
Xclkload71 clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload71/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload82 clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload82/Y sky130_fd_sc_hd__inv_6
XANTENNA_fanout1032_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload93 clknet_leaf_55_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload93/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_149_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09556__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10166__A1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09564__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout492_A net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08996_ _05056_ vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_145_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09308__B1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09861__A _05888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12698__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout757_A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09580__B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09617_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[2\]
+ net883 net869 net857 vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__and4_1
XFILLER_0_74_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08196__B team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[30\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout924_A net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1287_X net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12615__A0 _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09548_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[3\]
+ net660 net625 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[3\]
+ _05584_ vssd1 vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__a221o_1
XANTENNA__09087__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_120_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10626__C1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13830__B net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09479_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[4\]
+ net827 net803 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[4\]
+ _05515_ vssd1 vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout712_X net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13322__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11510_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[20\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[20\]
+ net1031 vssd1 vssd1 vccd1 vccd1 _07421_ sky130_fd_sc_hd__mux2_1
XANTENNA__11631__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14368__B1 _04082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12490_ net1660 _03612_ net211 vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11441_ net1 net1012 vssd1 vssd1 vccd1 vccd1 _07354_ sky130_fd_sc_hd__nor2_4
XFILLER_0_136_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14160_ _03963_ net907 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[9\]
+ sky130_fd_sc_hd__nor2_1
X_11372_ net957 _06756_ _06899_ _07309_ _06769_ vssd1 vssd1 vccd1 vccd1 _07310_ sky130_fd_sc_hd__o221a_1
XFILLER_0_34_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_104_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13111_ net270 net2671 net448 vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_169_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10323_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[24\] net904 _04238_
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[24\] _06344_ vssd1
+ vssd1 vccd1 vccd1 _06345_ sky130_fd_sc_hd__a221o_2
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14091_ _03957_ _03940_ vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__and2b_1
XFILLER_0_131_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_166_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_166_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09547__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input53_A wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13042_ net264 net2331 net456 vssd1 vssd1 vccd1 vccd1 _02600_ sky130_fd_sc_hd__mux2_1
X_10254_ _06124_ _06132_ net526 vssd1 vssd1 vccd1 vccd1 _06278_ sky130_fd_sc_hd__mux2_1
XANTENNA__13894__A2 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1201 net1202 vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__buf_2
X_17850_ clknet_leaf_98_wb_clk_i _03193_ _01546_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[32\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1212 net1213 vssd1 vssd1 vccd1 vccd1 net1212 sky130_fd_sc_hd__buf_4
X_10185_ _06003_ _06211_ vssd1 vssd1 vccd1 vccd1 _06212_ sky130_fd_sc_hd__or2_1
Xfanout1223 net1224 vssd1 vssd1 vccd1 vccd1 net1223 sky130_fd_sc_hd__buf_4
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1234 net1241 vssd1 vssd1 vccd1 vccd1 net1234 sky130_fd_sc_hd__clkbuf_4
X_16801_ clknet_leaf_148_wb_clk_i _02431_ _00497_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1245 net1252 vssd1 vssd1 vccd1 vccd1 net1245 sky130_fd_sc_hd__clkbuf_4
Xfanout1256 net1257 vssd1 vssd1 vccd1 vccd1 net1256 sky130_fd_sc_hd__buf_4
Xfanout1267 net1268 vssd1 vssd1 vccd1 vccd1 net1267 sky130_fd_sc_hd__buf_4
X_17781_ clknet_leaf_91_wb_clk_i _03124_ _01477_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1278 net1279 vssd1 vssd1 vccd1 vccd1 net1278 sky130_fd_sc_hd__clkbuf_2
X_14993_ net1189 vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__inv_2
Xfanout280 net281 vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__clkbuf_2
Xfanout291 net293 vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1289 net1291 vssd1 vssd1 vccd1 vccd1 net1289 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16732_ clknet_leaf_161_wb_clk_i _02362_ _00428_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12401__S _07852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13944_ _03805_ _03816_ _03817_ vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__and3_1
XANTENNA__08387__A net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13875_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[9\]
+ net559 net575 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[9\]
+ net986 vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__a221o_1
X_16663_ clknet_leaf_146_wb_clk_i _02293_ _00359_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_18402_ net915 vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__clkbuf_1
X_15614_ net1148 vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__inv_2
X_12826_ net324 net2783 net484 vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16594_ clknet_leaf_125_wb_clk_i _02224_ _00290_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09078__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18333_ net1322 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
XANTENNA__13740__B _06623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15545_ net1116 vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__inv_2
X_12757_ net321 net2634 net493 vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__mux2_1
XANTENNA__08825__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11541__A _07448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13232__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11708_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[9\] team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[10\]
+ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[14\] team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[6\]
+ vssd1 vssd1 vccd1 vccd1 _07520_ sky130_fd_sc_hd__or4b_1
X_15476_ net1172 vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__inv_2
X_18264_ clknet_leaf_38_wb_clk_i _03493_ _01959_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12688_ net2962 net340 vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17215_ clknet_leaf_152_wb_clk_i _02845_ _00911_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14427_ net1095 vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__inv_2
X_11639_ net25 net991 net918 net1923 vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__a22o_1
XANTENNA__14374__A3 _04146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18195_ clknet_leaf_33_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[16\]
+ _01890_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17146_ clknet_leaf_10_wb_clk_i _02776_ _00842_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_14358_ net375 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[7\]
+ _04096_ _04130_ _04111_ vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold706 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2120 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09250__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17585__D team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[22\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold717 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net2131 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13309_ net2272 net263 net428 vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__mux2_1
Xhold728 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2142 sky130_fd_sc_hd__dlygate4sd3_1
X_17077_ clknet_leaf_174_wb_clk_i _02707_ _00773_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold739 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[41\] vssd1 vssd1
+ vccd1 vccd1 net2153 sky130_fd_sc_hd__dlygate4sd3_1
X_14289_ _04062_ _06185_ _06108_ vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_55_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16028_ net1284 vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09002__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08850_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[18\]
+ net849 net798 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[18\]
+ _04907_ vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_51_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1406 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2820 sky130_fd_sc_hd__dlygate4sd3_1
X_08781_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[19\]
+ net643 net610 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__a22o_1
Xhold1417 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2831 sky130_fd_sc_hd__dlygate4sd3_1
X_17979_ clknet_leaf_106_wb_clk_i _03318_ _01675_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__dfrtp_1
Xhold1428 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net2842 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14299__A _04490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1439 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2853 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13407__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09402_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[6\]
+ net788 net769 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09069__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18288__1380 vssd1 vssd1 vccd1 vccd1 net1380 _18288__1380/LO sky130_fd_sc_hd__conb_1
X_09333_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[7\]
+ net705 net631 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08277__B1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[31\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_7_0_wb_clk_i_X clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08816__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_779 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13142__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09264_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[9\]
+ net824 net792 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[9\]
+ _05311_ vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08215_ _04232_ net962 _04271_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[15\]
+ _04155_ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__o311a_1
XANTENNA__18007__Q net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13022__A0 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09195_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[10\]
+ net668 net610 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__a22o_1
XANTENNA__12981__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout505_A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1247_A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08146_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[3\] team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[1\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[0\] vssd1 vssd1
+ vccd1 vccd1 _04229_ sky130_fd_sc_hd__and3b_1
XANTENNA__09856__A _04818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09241__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload160 clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload160/Y sky130_fd_sc_hd__inv_8
X_08077_ net1023 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__and2b_1
Xclkload171 clknet_leaf_89_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload171/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_141_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1035_X net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload182 clknet_leaf_91_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload182/Y sky130_fd_sc_hd__clkinv_2
Xclkload193 clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload193/Y sky130_fd_sc_hd__inv_8
XANTENNA__09529__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout495_X net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout874_A net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold11 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[26\]
+ vssd1 vssd1 vccd1 vccd1 net1425 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[28\]
+ vssd1 vssd1 vccd1 vccd1 net1436 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[12\]
+ vssd1 vssd1 vccd1 vccd1 net1447 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[8\] vssd1 vssd1
+ vccd1 vccd1 net1458 sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[15\]
+ net826 net741 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[15\]
+ _05040_ vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout662_X net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold55 team_05_WB.instance_to_wrap.BUSY_O vssd1 vssd1 vccd1 vccd1 net1469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[25\]
+ vssd1 vssd1 vccd1 vccd1 net1480 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13317__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold77 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[27\]
+ vssd1 vssd1 vccd1 vccd1 net1491 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ _07801_ _07798_ _07797_ vssd1 vssd1 vccd1 vccd1 _07802_ sky130_fd_sc_hd__nand3b_1
Xhold88 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[19\]
+ vssd1 vssd1 vccd1 vccd1 net1502 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1513 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09741__D net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10941_ _06364_ _06768_ _06898_ _06929_ net564 vssd1 vssd1 vccd1 vccd1 _06930_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout927_X net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13660_ net2263 net193 net385 vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10872_ _06805_ _06868_ _06802_ _06803_ vssd1 vssd1 vccd1 vccd1 _06869_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_156_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12611_ _07850_ _03672_ _07840_ vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__and3b_4
XFILLER_0_112_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13261__A0 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13591_ net2054 net306 net397 vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13052__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15330_ net1220 vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12542_ _07844_ _07849_ vssd1 vssd1 vccd1 vccd1 _03677_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09480__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15261_ net1087 vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__inv_2
X_12473_ net919 _07847_ vssd1 vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12891__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14212_ _04011_ net728 _04010_ vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__and3b_1
X_17000_ clknet_leaf_204_wb_clk_i _02630_ _00696_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11424_ net1753 _07314_ _07321_ vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__o21a_1
X_15192_ net1201 vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11575__B1 _07354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_8 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14143_ net1936 net503 net911 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[26\]
+ sky130_fd_sc_hd__and3_1
X_11355_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[3\] net508 _07297_
+ _07291_ vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08440__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10306_ net369 _06327_ _06325_ vssd1 vssd1 vccd1 vccd1 _06328_ sky130_fd_sc_hd__o21ai_2
X_14074_ _03940_ _03941_ vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__or2_1
X_11286_ net1844 net731 _07246_ vssd1 vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__o21a_1
XFILLER_0_120_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17902_ clknet_leaf_75_wb_clk_i _03245_ _01598_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13025_ net323 net2849 net460 vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__mux2_1
X_10237_ _06059_ _06261_ net531 vssd1 vssd1 vccd1 vccd1 _06262_ sky130_fd_sc_hd__mux2_1
Xfanout1020 net1021 vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__clkbuf_4
Xfanout1031 net1032 vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__clkbuf_4
Xfanout1042 net1047 vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__clkbuf_4
X_17833_ clknet_leaf_102_wb_clk_i _03176_ _01529_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[79\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13735__B _06706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1053 net1065 vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__buf_4
X_10168_ _06067_ _06070_ vssd1 vssd1 vccd1 vccd1 _06195_ sky130_fd_sc_hd__nor2_1
XFILLER_0_174_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1064 net1065 vssd1 vssd1 vccd1 vccd1 net1064 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13227__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1075 net1076 vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__clkbuf_4
Xfanout1086 net1107 vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12827__A0 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17764_ clknet_leaf_83_wb_clk_i _03107_ _01460_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1097 net1107 vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__clkbuf_4
X_14976_ net1197 vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__inv_2
XANTENNA__09299__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10099_ net349 net361 vssd1 vssd1 vccd1 vccd1 _06127_ sky130_fd_sc_hd__nand2_1
XANTENNA__09651__D net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_63_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16715_ clknet_leaf_188_wb_clk_i _02345_ _00411_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13927_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[6\] team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[5\]
+ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[7\] vssd1 vssd1 vccd1
+ vccd1 _03802_ sky130_fd_sc_hd__o21ai_1
X_17695_ clknet_leaf_86_wb_clk_i _03038_ _01391_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13751__A _05212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16646_ clknet_leaf_115_wb_clk_i _02276_ _00342_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13858_ net1563 net982 _03765_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[0\]
+ sky130_fd_sc_hd__o21a_1
X_12809_ net263 net2379 net484 vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16577_ clknet_leaf_150_wb_clk_i _02207_ _00273_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_146_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13789_ net1449 net974 net723 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[0\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_84_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14285__C _06464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18316_ net1408 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
XFILLER_0_32_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15528_ net1159 vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_79_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10158__Y _06185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18247_ clknet_leaf_38_wb_clk_i _03476_ _01942_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15459_ net1171 vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09759__B1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18178_ clknet_leaf_50_wb_clk_i net1048 _01873_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09223__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold503 net82 vssd1 vssd1 vccd1 vccd1 net1917 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold514 net99 vssd1 vssd1 vccd1 vccd1 net1928 sky130_fd_sc_hd__dlygate4sd3_1
X_17129_ clknet_leaf_20_wb_clk_i _02759_ _00825_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold525 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[13\] vssd1
+ vssd1 vccd1 vccd1 net1939 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold536 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net1950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 _03302_ vssd1 vssd1 vccd1 vccd1 net1961 sky130_fd_sc_hd__dlygate4sd3_1
X_09951_ _05977_ _05978_ _05979_ vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__nor3_1
Xhold558 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 net1972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 net1983 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11318__B1 _07127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08902_ _04966_ _04944_ vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__and2b_2
XTAP_TAPCELL_ROW_70_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09882_ _04594_ _05910_ vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__nand2_1
X_08833_ _04359_ _04901_ vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__nand2_1
Xhold1203 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1214 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1225 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net2639 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout288_A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13137__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1236 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2650 sky130_fd_sc_hd__dlygate4sd3_1
X_08764_ _04832_ _04834_ _04835_ vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__or3_1
Xhold1247 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1258 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1269 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 net2683 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08498__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12976__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08695_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[22\]
+ net678 net669 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout455_A _03713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_146_Right_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09203__X _05256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout622_A net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09316_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[8\]
+ net776 net758 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__a22o_1
XFILLER_0_165_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09247_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[9\]
+ net666 net603 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08670__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout410_X net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14492__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13600__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09178_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[11\]
+ net752 net733 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[11\]
+ _05218_ vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__a221o_1
XANTENNA__09214__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08129_ _04214_ net154 net153 vssd1 vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__or3b_2
XANTENNA__08422__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10525__A _04265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11140_ _07087_ _07079_ _07075_ vssd1 vssd1 vccd1 vccd1 _07106_ sky130_fd_sc_hd__and3b_4
XANTENNA__11309__B1 _07130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__clkbuf_4
X_11071_ _07036_ _07037_ vssd1 vssd1 vccd1 vccd1 _07038_ sky130_fd_sc_hd__and2_2
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__clkbuf_4
XANTENNA__08725__A1 _04344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10022_ _04157_ _05923_ vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__nor2_4
XANTENNA__09752__C net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13047__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14830_ net1187 vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input16_A DAT_I[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11973_ _07766_ _07780_ _07782_ _07784_ vssd1 vssd1 vccd1 vccd1 _07785_ sky130_fd_sc_hd__and4_1
XANTENNA__12886__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14761_ net1221 vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__inv_2
XANTENNA__08489__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13482__A0 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16500_ clknet_leaf_112_wb_clk_i _02130_ _00196_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_13712_ net900 _06557_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[12\]
+ sky130_fd_sc_hd__nor2_1
X_10924_ _06273_ _06915_ net957 vssd1 vssd1 vccd1 vccd1 _06916_ sky130_fd_sc_hd__mux2_1
X_17480_ clknet_leaf_37_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[15\]
+ _01176_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_14692_ net1236 vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16431_ clknet_leaf_137_wb_clk_i _02061_ _00127_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10855_ _06829_ _06851_ _06828_ vssd1 vssd1 vccd1 vccd1 _06852_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_67_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13643_ net2889 net275 net391 vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16362_ clknet_leaf_17_wb_clk_i _01992_ _00058_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13574_ net2134 net260 net397 vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__mux2_1
X_10786_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[27\] net1041 vssd1
+ vssd1 vccd1 vccd1 _06783_ sky130_fd_sc_hd__and2_1
XANTENNA__10599__A1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09453__A2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18101_ clknet_leaf_52_wb_clk_i _03424_ _01797_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[18\]
+ sky130_fd_sc_hd__dfrtp_2
X_12525_ net1763 _03632_ net208 vssd1 vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__mux2_1
XANTENNA__15498__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15313_ net1216 vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__inv_2
X_16293_ net1154 vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__inv_2
XANTENNA__11260__A2 _07103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12474__X _03673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_181_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_181_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_81_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13510__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18032_ clknet_leaf_97_wb_clk_i _03371_ _01728_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12456_ net1665 _03632_ net212 vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__mux2_1
X_15244_ net1072 vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_110_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_110_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11407_ _07329_ net1966 vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15175_ net1199 vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__inv_2
XANTENNA__08413__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12387_ net1631 _03663_ _07852_ vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12353__C _03645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09646__D net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14126_ _03798_ _03989_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[12\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_91_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11338_ team_05_WB.instance_to_wrap.total_design.keypad0.next_rows\[1\] team_05_WB.instance_to_wrap.total_design.keypad0.next_rows\[3\]
+ team_05_WB.instance_to_wrap.total_design.keypad0.next_rows\[2\] vssd1 vssd1 vccd1
+ vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.next_rows\[0\] sky130_fd_sc_hd__nand3_1
XFILLER_0_10_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13746__A _05213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14057_ _03924_ _03925_ vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__nand2_1
X_11269_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[2\] _07092_ _07101_
+ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[10\] vssd1 vssd1 vccd1
+ vccd1 _07230_ sky130_fd_sc_hd__a22o_1
XFILLER_0_158_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13008_ net258 net2433 net460 vssd1 vssd1 vccd1 vccd1 _02633_ sky130_fd_sc_hd__mux2_1
XANTENNA__11537__Y _07448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10523__B2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[14\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17816_ clknet_leaf_90_wb_clk_i _03159_ _01512_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[126\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17747_ clknet_leaf_90_wb_clk_i _03090_ _01443_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12796__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14959_ net1282 vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__inv_2
X_08480_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[27\]
+ net603 net595 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__a22o_1
X_17678_ clknet_leaf_84_wb_clk_i _03021_ _01374_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[116\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16629_ clknet_leaf_22_wb_clk_i _02259_ _00325_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1068 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_28_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09101_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[12\]
+ net643 net611 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_135_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11251__A2 _07117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08652__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13420__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09032_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[14\]
+ net770 net743 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold300 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[21\] vssd1 vssd1
+ vccd1 vccd1 net1714 sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 team_05_WB.instance_to_wrap.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 net1725
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout203_A net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold322 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[29\] vssd1 vssd1
+ vccd1 vccd1 net1736 sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[58\] vssd1 vssd1
+ vccd1 vccd1 net1747 sky130_fd_sc_hd__dlygate4sd3_1
Xhold344 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[51\] vssd1 vssd1
+ vccd1 vccd1 net1758 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[5\] vssd1 vssd1
+ vccd1 vccd1 net1769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 net89 vssd1 vssd1 vccd1 vccd1 net1780 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold377 team_05_WB.instance_to_wrap.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 net1791
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold388 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[92\] vssd1 vssd1
+ vccd1 vccd1 net1802 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout802 net805 vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__buf_4
Xhold399 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[75\] vssd1 vssd1
+ vccd1 vccd1 net1813 sky130_fd_sc_hd__dlygate4sd3_1
X_09934_ _05831_ _05962_ _05832_ vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__o21ai_1
Xfanout813 _04390_ vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__buf_4
XANTENNA__16032__A net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout824 net825 vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_37_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout835 net836 vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__clkbuf_4
Xfanout846 _04373_ vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__clkbuf_4
X_09865_ _05888_ _05893_ _05892_ _04757_ vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__a211o_1
Xfanout857 net859 vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__buf_2
XANTENNA_input8_A DAT_I[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09572__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1000 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2414 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout572_A net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout868 _04289_ vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__buf_2
Xhold1011 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2425 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout879 net882 vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__buf_2
Xhold1022 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2436 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1033 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2447 sky130_fd_sc_hd__dlygate4sd3_1
X_08816_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[18\]
+ net695 net632 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[18\]
+ _04882_ vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__a221o_1
X_09796_ _05826_ vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__inv_2
Xhold1044 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 net2458 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1055 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net2469 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1066 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1077 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2491 sky130_fd_sc_hd__dlygate4sd3_1
X_08747_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[21\]
+ net819 net807 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__a22o_1
Xhold1088 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2502 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1099 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net2513 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout837_A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout458_X net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1081 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08678_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[23\]
+ net835 _04751_ net855 vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_159_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1054 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout625_X net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08891__B1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_46_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10640_ _06010_ _06022_ vssd1 vssd1 vccd1 vccd1 _06645_ sky130_fd_sc_hd__nand2_1
XANTENNA__09435__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1030 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11242__A2 _07100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10571_ _06018_ _06029_ vssd1 vssd1 vccd1 vccd1 _06580_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12310_ _07894_ _08022_ _03537_ _03603_ vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__o22a_4
XANTENNA__13330__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13290_ net330 net2840 net434 vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__mux2_1
XANTENNA__09747__C net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12241_ _03512_ _03533_ _03535_ _03532_ vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_31_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12172_ _07968_ _07972_ vssd1 vssd1 vccd1 vccd1 _07984_ sky130_fd_sc_hd__and2b_1
XFILLER_0_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11123_ net1934 _07031_ _07086_ _07089_ vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_55_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16980_ clknet_leaf_119_wb_clk_i _02610_ _00676_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11054_ net957 _06729_ _07021_ vssd1 vssd1 vccd1 vccd1 _07022_ sky130_fd_sc_hd__o21ai_1
X_15931_ net1301 vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__inv_2
X_10005_ net377 net367 vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__nand2_1
X_15862_ net1267 vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__inv_2
XANTENNA__08947__X team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[16\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17601_ clknet_leaf_79_wb_clk_i _02972_ _01297_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_14813_ net1088 vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__inv_2
X_15793_ net1276 vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__inv_2
XANTENNA__10269__B1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13505__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17532_ clknet_leaf_81_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[3\]
+ _01228_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14744_ net1244 vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__inv_2
X_11956_ _07527_ _07761_ vssd1 vssd1 vccd1 vccd1 _07768_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_28_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13207__A0 _06461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17463_ clknet_leaf_58_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[31\]
+ _01159_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10907_ net963 _06185_ _06901_ vssd1 vssd1 vccd1 vccd1 _06902_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14675_ net1215 vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__inv_2
XANTENNA__08882__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11887_ _07669_ _07671_ _07664_ vssd1 vssd1 vccd1 vccd1 _07699_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_168_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16414_ clknet_leaf_163_wb_clk_i _02044_ _00110_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10838_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[3\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06835_ sky130_fd_sc_hd__nand2_1
X_13626_ net2082 net200 net390 vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17394_ clknet_leaf_65_wb_clk_i net1425 _01090_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09426__A2 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11233__A2 _07116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16345_ clknet_leaf_10_wb_clk_i _01975_ _00041_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13557_ net1946 net326 net401 vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__mux2_1
X_10769_ net383 _06766_ vssd1 vssd1 vccd1 vccd1 _06767_ sky130_fd_sc_hd__and2_1
XFILLER_0_109_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13240__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10441__B1 _04275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12508_ _07840_ _07843_ vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__nand2_8
XFILLER_0_70_836 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16276_ net1147 vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__inv_2
X_13488_ net331 net2469 net410 vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__mux2_1
X_18015_ clknet_leaf_64_wb_clk_i _03354_ _01711_ vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__dfrtp_1
X_12439_ _07840_ _07850_ _03669_ vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__and3_4
XFILLER_0_113_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15227_ net1099 vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_130_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14860__A net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15158_ net1101 vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__inv_2
XANTENNA__17593__D team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[30\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14109_ _03949_ _03973_ _03972_ vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15089_ net1188 vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__inv_2
XANTENNA__12497__A1 _07798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11708__B team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[10\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08289__B team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[22\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09650_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[1\]
+ net946 net1013 net927 vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__and4_1
X_08601_ _04675_ vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__inv_2
XANTENNA__13923__B _07451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09581_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[2\]
+ net950 net936 net929 vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__and4_1
X_18397__1371 vssd1 vssd1 vccd1 vccd1 _18397__1371/HI net1371 sky130_fd_sc_hd__conb_1
XANTENNA__13415__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08532_ _04602_ _04604_ _04606_ _04608_ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_26_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08463_ _04535_ _04537_ _04539_ _04541_ vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__or4_2
XANTENNA__08873__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08394_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[29\]
+ net669 net631 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[29\]
+ _04473_ vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__a221o_1
XANTENNA__09417__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08625__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout320_A _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13150__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1062_A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout418_A net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10346__Y _06367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09567__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09015_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[14\]
+ net667 net622 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[14\]
+ _05062_ vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__a221o_1
XFILLER_0_171_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold130 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[6\] vssd1 vssd1
+ vccd1 vccd1 net1544 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold141 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[28\]
+ vssd1 vssd1 vccd1 vccd1 net1555 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_37_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_112_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09050__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold152 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[11\]
+ vssd1 vssd1 vccd1 vccd1 net1566 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 team_05_WB.instance_to_wrap.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 net1577
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout787_A _04400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold174 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[28\] vssd1 vssd1
+ vccd1 vccd1 net1588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[0\] vssd1
+ vssd1 vccd1 vccd1 net1599 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09583__B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold196 team_05_WB.instance_to_wrap.total_design.core.data_access vssd1 vssd1 vccd1
+ vccd1 net1610 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13817__C net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout610 _04319_ vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__buf_6
Xfanout621 net624 vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__clkbuf_8
Xfanout632 net633 vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__clkbuf_8
X_09917_ _05735_ _05944_ _05945_ vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__a21o_1
Xfanout643 _04311_ vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_109_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout654 net655 vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_109_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09353__A1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[27\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout665 _04305_ vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12440__D _03659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout676 net679 vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__buf_6
X_09848_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[20\]
+ net590 _05869_ _05878_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[20\]
+ sky130_fd_sc_hd__o22a_4
Xfanout687 net690 vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__clkbuf_8
Xfanout698 _04295_ vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_126_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout742_X net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13833__B net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09779_ _05442_ _05463_ vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__and2b_1
XFILLER_0_38_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11634__A team_05_WB.instance_to_wrap.wishbone.curr_state\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13325__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11810_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[5\] net997 vssd1
+ vssd1 vccd1 vccd1 _07622_ sky130_fd_sc_hd__nand2_1
X_12790_ net323 net1963 net489 vssd1 vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09656__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11741_ net550 _07552_ vssd1 vssd1 vccd1 vccd1 _07553_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_1_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08864__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10671__B1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11672_ team_05_WB.EN_VAL_REG net1049 net507 _07486_ vssd1 vssd1 vccd1 vccd1 _07487_
+ sky130_fd_sc_hd__nand4_1
X_14460_ net1074 vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__inv_2
XANTENNA__09408__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13411_ net2743 net271 net416 vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__mux2_1
X_10623_ _06560_ _06628_ net529 vssd1 vssd1 vccd1 vccd1 _06629_ sky130_fd_sc_hd__mux2_1
X_14391_ net1545 vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11215__A2 _07099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_76_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13060__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16130_ net1303 vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__inv_2
X_13342_ net263 net2877 net424 vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10554_ _06412_ net332 _06561_ net335 vssd1 vssd1 vccd1 vccd1 _06564_ sky130_fd_sc_hd__o22a_1
XFILLER_0_51_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16061_ net1262 vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__inv_2
X_13273_ net247 net2651 net434 vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10485_ _06494_ _06498_ net382 vssd1 vssd1 vccd1 vccd1 _06499_ sky130_fd_sc_hd__o21a_2
XFILLER_0_106_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12224_ _08015_ _08019_ vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15012_ net1230 vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09041__B1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[14\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08395__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12155_ _07963_ _07966_ vssd1 vssd1 vccd1 vccd1 _07967_ sky130_fd_sc_hd__nand2_1
X_11106_ _07052_ _07058_ vssd1 vssd1 vccd1 vccd1 _07073_ sky130_fd_sc_hd__and2b_2
XANTENNA__11528__B _07434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12479__A1 _03651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16963_ clknet_leaf_198_wb_clk_i _02593_ _00659_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_12086_ _07892_ _07894_ _07896_ vssd1 vssd1 vccd1 vccd1 _07898_ sky130_fd_sc_hd__or3_1
XFILLER_0_21_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11037_ net1046 _06686_ _07007_ net959 vssd1 vssd1 vccd1 vccd1 _07008_ sky130_fd_sc_hd__o211a_1
X_15914_ net1288 vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16894_ clknet_leaf_184_wb_clk_i _02524_ _00590_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08552__C1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13743__B _06572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15845_ net1270 vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13235__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15016__A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15776_ net1275 vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12988_ net319 net2409 net466 vssd1 vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__mux2_1
XANTENNA__12100__B1 _07864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17515_ clknet_leaf_73_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[18\]
+ _01211_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[18\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_82_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14727_ net1176 vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__inv_2
X_11939_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[1\] net999 vssd1
+ vssd1 vccd1 vccd1 _07751_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12651__B2 _07351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17446_ clknet_leaf_60_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[14\]
+ _01142_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10662__B1 _06055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14658_ net1217 vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_60_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17588__D team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[25\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09301__X _05350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12403__A1 _03623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11206__A2 _07092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13609_ net2773 net271 net392 vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17377_ clknet_leaf_81_wb_clk_i net1427 _01073_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08607__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14589_ net1089 vssd1 vssd1 vccd1 vccd1 _00219_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16328_ net1126 vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09280__B1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08291__C net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16259_ net1119 vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wire376_X net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09032__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08386__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[30\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11438__B net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09702_ net512 _05731_ vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_156_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09633_ net527 net523 vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_104_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13145__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09564_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[2\]
+ net944 net939 _04418_ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__and4_1
XANTENNA__09099__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_8__f_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08515_ net570 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[27\]
+ _04362_ vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__o21a_1
XFILLER_0_66_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_110_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12642__A1 _07836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09495_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[4\]
+ net684 net622 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__a22o_1
XANTENNA__08846__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12984__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1277_A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08310__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10653__B1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08446_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[28\]
+ net693 net685 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_173_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08377_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[30\]
+ net847 net823 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[30\]
+ _04457_ vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__a221o_1
XANTENNA__09578__B net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout702_A _04293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout323_X net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1065_X net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09271__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10270_ _06289_ _06293_ _04265_ vssd1 vssd1 vccd1 vccd1 _06294_ sky130_fd_sc_hd__o21a_2
XANTENNA__09023__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout692_X net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08377__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09744__D net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout440 _03716_ vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__buf_8
Xfanout451 _03714_ vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__buf_4
Xfanout462 _03711_ vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__buf_6
X_13960_ _03831_ _03832_ vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__or2_1
Xfanout473 _03706_ vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__clkbuf_4
Xfanout484 _03703_ vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_6_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08534__C1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout495 _03699_ vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__buf_4
X_12911_ net271 net2940 net472 vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__mux2_1
X_13891_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[17\]
+ net558 net574 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[17\]
+ net985 vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__a221o_1
XANTENNA__13055__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15630_ net1246 vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__inv_2
XANTENNA__10892__B1 _04170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12842_ net264 net2313 net480 vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__mux2_1
XANTENNA__09629__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15561_ net1118 vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__inv_2
X_12773_ net255 net2814 net488 vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__mux2_1
XANTENNA__08837__B1 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17300_ clknet_leaf_128_wb_clk_i _02930_ _00996_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_14512_ net1092 vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__inv_2
X_18280_ net107 vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__clkbuf_1
X_11724_ _07535_ vssd1 vssd1 vccd1 vccd1 _07536_ sky130_fd_sc_hd__inv_2
X_15492_ net1158 vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_199_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17231_ clknet_leaf_141_wb_clk_i _02861_ _00927_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_11655_ net7 net991 net918 net1906 vssd1 vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__a22o_1
X_14443_ net1068 vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__inv_2
XANTENNA__10708__A net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_88_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_142_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17162_ clknet_leaf_195_wb_clk_i _02792_ _00858_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10606_ _06544_ _06612_ net529 vssd1 vssd1 vccd1 vccd1 _06613_ sky130_fd_sc_hd__mux2_1
X_11586_ net1977 net1006 _07367_ net357 vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__a22o_1
X_14374_ net1022 _04268_ _04146_ _04247_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.branch_ff
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09262__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16113_ net1135 vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__inv_2
X_10537_ _05833_ _06056_ _06198_ _06509_ _06547_ vssd1 vssd1 vccd1 vccd1 _06548_ sky130_fd_sc_hd__a221o_1
XFILLER_0_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_17_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13325_ net2785 net322 net431 vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__mux2_1
X_17093_ clknet_leaf_175_wb_clk_i _02723_ _00789_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16044_ net1287 vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__inv_2
X_13256_ net315 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[5\]
+ net439 vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__mux2_1
XANTENNA__09014__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10468_ _05014_ _05966_ _05968_ vssd1 vssd1 vccd1 vccd1 _06482_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08368__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12207_ _08014_ _08018_ _08012_ vssd1 vssd1 vccd1 vccd1 _08019_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_36_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13187_ net315 net2830 net443 vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10399_ net348 _06413_ _06416_ vssd1 vssd1 vccd1 vccd1 _06417_ sky130_fd_sc_hd__o21ai_1
X_12138_ _07943_ _07949_ _07947_ vssd1 vssd1 vccd1 vccd1 _07950_ sky130_fd_sc_hd__o21ai_2
X_17995_ clknet_leaf_82_wb_clk_i _03334_ _01691_ vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13754__A _05212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09951__B _05978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12069_ _07868_ _07879_ vssd1 vssd1 vccd1 vccd1 _07881_ sky130_fd_sc_hd__or2_1
X_16946_ clknet_leaf_120_wb_clk_i _02576_ _00642_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14310__B2 _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16877_ clknet_leaf_160_wb_clk_i _02507_ _00573_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09670__C net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08540__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15828_ net1307 vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__inv_2
X_15759_ net1299 vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__inv_2
XANTENNA__08828__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12657__X _03693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08300_ net942 net930 net925 vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__and3_1
X_09280_ net572 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[9\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[9\] vssd1 vssd1 vccd1
+ vccd1 _05329_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08231_ net878 net864 net860 vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__and3_4
X_17429_ clknet_leaf_60_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[29\]
+ _01125_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_166_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08162_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[3\] team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[1\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[0\] _04242_ vssd1
+ vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__and4_1
XFILLER_0_28_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08093_ net1023 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__and2b_1
XFILLER_0_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16305__A net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_11__f_wb_clk_i_X clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkload50 clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload50/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_77_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09005__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload61 clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload61/Y sky130_fd_sc_hd__inv_16
Xclkload72 clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload72/Y sky130_fd_sc_hd__clkinv_2
Xclkload83 clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload83/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload94 clknet_leaf_56_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload94/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__08359__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10353__A _06051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12560__A0 _03632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09564__D _04418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12979__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08995_ _05034_ _05055_ vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_10_Left_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout485_A _03703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09580__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout652_A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08531__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09616_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[2\]
+ net876 net867 net860 vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__and4_1
XFILLER_0_92_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09547_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[3\]
+ net652 net648 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__a22o_1
XANTENNA__08819__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout440_X net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout538_X net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13603__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09492__B1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09478_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[4\]
+ net796 net739 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08429_ _04504_ _04505_ _04506_ _04508_ vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout705_X net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11440_ _07349_ _07351_ team_05_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 _07353_ sky130_fd_sc_hd__o21ai_2
Xclkload0 clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload0/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09244__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11371_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[0\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[0\]
+ vssd1 vssd1 vccd1 vccd1 _07309_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16215__A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10322_ net895 _06343_ vssd1 vssd1 vccd1 vccd1 _06344_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13110_ net267 net2892 net448 vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__mux2_1
X_14090_ _03938_ _03954_ _03955_ _03953_ vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__a211o_1
XANTENNA__09755__C net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13041_ net257 net2333 net457 vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__mux2_1
X_10253_ net526 _06116_ vssd1 vssd1 vccd1 vccd1 _06277_ sky130_fd_sc_hd__nand2_1
XANTENNA__12551__A0 _03657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input46_A wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10184_ _06207_ _06210_ net372 vssd1 vssd1 vccd1 vccd1 _06211_ sky130_fd_sc_hd__mux2_1
Xfanout1202 net1211 vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__clkbuf_2
Xfanout1213 net1241 vssd1 vssd1 vccd1 vccd1 net1213 sky130_fd_sc_hd__buf_4
XANTENNA__12889__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1224 net1225 vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__buf_4
Xfanout1235 net1237 vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__buf_4
X_16800_ clknet_leaf_128_wb_clk_i _02430_ _00496_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08770__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1246 net1247 vssd1 vssd1 vccd1 vccd1 net1246 sky130_fd_sc_hd__buf_4
X_17780_ clknet_leaf_84_wb_clk_i _03123_ _01476_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09771__B _05801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1257 net1279 vssd1 vssd1 vccd1 vccd1 net1257 sky130_fd_sc_hd__buf_4
X_14992_ net1092 vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_135_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_135_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout1268 net1271 vssd1 vssd1 vccd1 vccd1 net1268 sky130_fd_sc_hd__clkbuf_2
Xfanout270 net273 vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_31_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1279 net1312 vssd1 vssd1 vccd1 vccd1 net1279 sky130_fd_sc_hd__buf_2
Xfanout281 _06571_ vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout292 net293 vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__clkbuf_2
X_16731_ clknet_leaf_190_wb_clk_i _02361_ _00427_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13943_ _03811_ _03815_ vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__nand2_1
XANTENNA__08522__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16662_ clknet_leaf_139_wb_clk_i _02292_ _00358_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13874_ net1463 net983 _03773_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[8\]
+ sky130_fd_sc_hd__o21a_1
X_18401_ net914 vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_1
X_15613_ net1149 vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__inv_2
XANTENNA__12606__A1 _07816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12825_ net321 net2968 net484 vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__mux2_1
X_16593_ clknet_leaf_121_wb_clk_i _02223_ _00289_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13513__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18332_ net1321 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
X_15544_ net1132 vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12756_ net311 net2116 net492 vssd1 vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__mux2_1
XANTENNA__09483__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17489__Q team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[24\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_7__f_wb_clk_i_X clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_45_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11290__B1 _07128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11541__B _07451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11707_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[11\] _07379_ _07447_
+ _07478_ vssd1 vssd1 vccd1 vccd1 _07519_ sky130_fd_sc_hd__or4_2
X_18263_ clknet_leaf_37_wb_clk_i _03492_ _01958_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[17\]
+ sky130_fd_sc_hd__dfrtp_4
X_15475_ net1172 vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12687_ net2490 net340 vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__and2_1
XANTENNA__09649__D net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17214_ clknet_leaf_163_wb_clk_i _02844_ _00910_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_14426_ net1062 vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__inv_2
X_11638_ net26 net990 net917 net1609 vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__o22a_1
X_18194_ clknet_leaf_37_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[15\]
+ _01889_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09235__B1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08589__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13749__A _05212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17145_ clknet_leaf_9_wb_clk_i _02775_ _00841_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14357_ _04100_ _04114_ _04129_ _04102_ _04097_ vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__o221a_1
X_11569_ net1922 net1004 net727 _07414_ vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12790__A0 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold707 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 net2121 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11593__B2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[31\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13308_ net2476 net255 net428 vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold718 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net2132 sky130_fd_sc_hd__dlygate4sd3_1
Xhold729 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 net2143 sky130_fd_sc_hd__dlygate4sd3_1
X_17076_ clknet_leaf_128_wb_clk_i _02706_ _00772_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_14288_ _06219_ _06273_ _04052_ _04061_ vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__or4_1
XFILLER_0_126_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16027_ net1284 vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__inv_2
X_13239_ net226 net2165 net437 vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12799__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11556__X _07467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08761__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08780_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[19\]
+ net691 net675 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[19\]
+ _04850_ vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__a221o_1
Xhold1407 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2821 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17978_ clknet_leaf_106_wb_clk_i _03317_ _01674_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__dfrtp_1
Xhold1418 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2832 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1429 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2843 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14295__B1 _04656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14299__B _04510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16929_ clknet_leaf_151_wb_clk_i _02559_ _00625_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11648__A2 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10620__B _06328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08513__A2 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_140_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09401_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[6\]
+ net813 net755 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__a22o_1
XFILLER_0_172_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10608__B1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11732__A team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[11\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13423__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09332_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[7\]
+ net680 net638 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05379_ sky130_fd_sc_hd__a22o_1
XANTENNA__09474__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11281__B1 _07111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09263_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[9\]
+ net747 net742 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[9\]
+ _05312_ vssd1 vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout233_A _06367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08214_ net885 net868 net861 vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09194_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[10\]
+ net682 net597 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[10\]
+ _05246_ vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__a221o_1
XFILLER_0_145_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08145_ _04228_ _04218_ net2957 vssd1 vssd1 vccd1 vccd1 _03471_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout400_A net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1142_A net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16035__A net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08076_ net1025 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[23\]
+ net971 _04187_ vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__a22o_1
Xclkload150 clknet_leaf_135_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload150/Y sky130_fd_sc_hd__bufinv_16
Xclkload161 clknet_leaf_77_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload161/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__09575__C net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload172 clknet_leaf_90_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload172/X sky130_fd_sc_hd__clkbuf_8
Xclkload183 clknet_leaf_92_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload183/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_101_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09872__A _04656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_164_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout390_X net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout867_A net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout488_X net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[30\]
+ vssd1 vssd1 vccd1 vccd1 net1426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[11\]
+ vssd1 vssd1 vccd1 vccd1 net1437 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12502__S _03673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold34 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[20\]
+ vssd1 vssd1 vccd1 vccd1 net1448 sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[15\]
+ net806 net794 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05040_ sky130_fd_sc_hd__a22o_1
Xhold45 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[31\]
+ vssd1 vssd1 vccd1 vccd1 net1459 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[10\] vssd1 vssd1
+ vccd1 vccd1 net1470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[12\] vssd1 vssd1
+ vccd1 vccd1 net1481 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11639__A2 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold78 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[27\]
+ vssd1 vssd1 vccd1 vccd1 net1492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[3\]
+ vssd1 vssd1 vccd1 vccd1 net1503 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout655_X net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08504__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10940_ _06876_ _06928_ vssd1 vssd1 vccd1 vccd1 _06929_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10871_ _06804_ _06867_ vssd1 vssd1 vccd1 vccd1 _06868_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout822_X net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13333__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12610_ _03623_ net1855 net203 vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__mux2_1
XANTENNA__15114__A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13590_ net2736 net324 net397 vssd1 vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10529__Y _06540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11272__B1 _07097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12541_ net1638 _03623_ net208 vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15260_ net1083 vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12472_ net1634 _03623_ net212 vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14211_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[11\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[10\]
+ _04008_ vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__and3_1
XFILLER_0_163_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11423_ _07322_ _07340_ vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__nor2_1
X_15191_ net1102 vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_9 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11354_ _07289_ team_05_WB.instance_to_wrap.total_design.keypad0.next_rows\[3\] net508
+ vssd1 vssd1 vccd1 vccd1 _07297_ sky130_fd_sc_hd__a21oi_1
X_14142_ net1725 net503 net911 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[25\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_105_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10305_ net525 _06226_ _06326_ vssd1 vssd1 vccd1 vccd1 _06327_ sky130_fd_sc_hd__o21a_1
XFILLER_0_120_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08991__A2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11285_ _07234_ _07240_ _07241_ _07245_ vssd1 vssd1 vccd1 vccd1 _07246_ sky130_fd_sc_hd__or4_1
X_14073_ _03938_ _03939_ _03914_ _03918_ vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__a211oi_1
XANTENNA__12760__X _03700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17901_ clknet_leaf_102_wb_clk_i _03244_ _01597_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10236_ _06260_ vssd1 vssd1 vccd1 vccd1 _06261_ sky130_fd_sc_hd__inv_2
X_13024_ net309 net2921 net460 vssd1 vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__mux2_1
XANTENNA__10535__C1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1010 net1011 vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__clkbuf_2
Xfanout1021 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[12\] vssd1
+ vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__clkbuf_4
X_17832_ clknet_leaf_92_wb_clk_i _03175_ _01528_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[78\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08743__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13508__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1032 net1036 vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__buf_2
XANTENNA__12412__S net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10167_ _04513_ _04514_ net510 _06193_ vssd1 vssd1 vccd1 vccd1 _06194_ sky130_fd_sc_hd__o31a_1
Xfanout1043 net1047 vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__clkbuf_2
Xfanout1054 net1055 vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__buf_4
Xfanout1065 net1108 vssd1 vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__buf_2
X_17763_ clknet_leaf_77_wb_clk_i _03106_ _01459_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1076 net1078 vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__buf_2
Xfanout1087 net1094 vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__buf_4
X_14975_ net1179 vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__inv_2
X_10098_ _05256_ net361 vssd1 vssd1 vccd1 vccd1 _06126_ sky130_fd_sc_hd__or2_1
Xfanout1098 net1100 vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__buf_4
X_16714_ clknet_leaf_195_wb_clk_i _02344_ _00410_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13926_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[10\] net979 team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__o21a_1
X_17694_ clknet_leaf_87_wb_clk_i _03037_ _01390_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[68\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13751__B _06424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16645_ clknet_leaf_180_wb_clk_i _02275_ _00341_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13857_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[0\]
+ net560 net576 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[0\]
+ net987 vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__a221o_1
XANTENNA__12648__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13243__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12808_ net255 net2417 net484 vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16576_ clknet_leaf_132_wb_clk_i _02206_ _00272_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09456__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13788_ _03760_ _03748_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.next_write
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_8_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18315_ net1407 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
X_15527_ net1159 vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__inv_2
XANTENNA__11263__B1 _07130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12739_ net254 net2689 net492 vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_32_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_32_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14863__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18246_ clknet_leaf_36_wb_clk_i _03475_ _01941_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_44_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15458_ net1171 vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14409_ net953 _04360_ _04346_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[22\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18177_ clknet_leaf_50_wb_clk_i net1535 _01872_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15389_ net1092 vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold504 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[13\] vssd1 vssd1
+ vccd1 vccd1 net1918 sky130_fd_sc_hd__dlygate4sd3_1
X_17128_ clknet_leaf_204_wb_clk_i _02758_ _00824_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold515 team_05_WB.instance_to_wrap.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 net1929
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold526 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1940 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold537 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net1951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1962 sky130_fd_sc_hd__dlygate4sd3_1
X_09950_ _04818_ _04838_ vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__and2b_1
XANTENNA__08982__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17059_ clknet_leaf_199_wb_clk_i _02689_ _00755_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold559 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net1973 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12515__A0 _07791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08901_ net571 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[17\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[17\] vssd1 vssd1 vccd1
+ vccd1 _04966_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_70_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ _04573_ _04593_ vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_70_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08734__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13418__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08832_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[18\] _04357_
+ vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1204 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2618 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1215 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 net2629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1226 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 net2640 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1237 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2651 sky130_fd_sc_hd__dlygate4sd3_1
X_08763_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[21\]
+ net757 net753 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[21\]
+ _04820_ vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__a221o_1
Xhold1248 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2662 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10350__B _06369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1259 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 net2673 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08694_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[22\]
+ net619 net615 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[22\]
+ _04766_ vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__a221o_1
XFILLER_0_164_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_68_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout350_A _03717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1092_A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13153__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout448_A _03714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09447__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10349__Y _06369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11254__B1 _07116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09315_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[8\]
+ net839 net773 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[8\]
+ _05362_ vssd1 vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12992__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout615_A _04318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09867__A net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09246_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[9\]
+ net688 net657 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[9\]
+ _05296_ vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__a221o_1
XFILLER_0_133_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09177_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[11\]
+ net849 net845 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[11\]
+ _05220_ vssd1 vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__a221o_1
XANTENNA__09586__B net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout403_X net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08128_ net154 net153 net152 net151 vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__and4b_1
XFILLER_0_102_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10765__C1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10525__B _06536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08059_ net1027 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout1312_X net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11070_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[3\] _07035_
+ vssd1 vssd1 vccd1 vccd1 _07037_ sky130_fd_sc_hd__or2_2
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout772_X net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10021_ net369 _06048_ vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__nand2_1
XANTENNA__08725__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[22\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10541__A net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09752__D net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14760_ net1218 vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11972_ _07728_ _07743_ _07783_ net343 vssd1 vssd1 vccd1 vccd1 _07784_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_99_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13711_ net901 _06572_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[11\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__09150__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10923_ net1044 _06880_ _06913_ _06914_ vssd1 vssd1 vccd1 vccd1 _06915_ sky130_fd_sc_hd__a31o_1
XFILLER_0_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14691_ net1207 vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13063__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16430_ clknet_leaf_170_wb_clk_i _02060_ _00126_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13642_ net2574 net273 net388 vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__mux2_1
X_10854_ _06831_ _06850_ _06830_ vssd1 vssd1 vccd1 vccd1 _06851_ sky130_fd_sc_hd__a21bo_1
XANTENNA__09438__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16361_ clknet_leaf_16_wb_clk_i _01991_ _00057_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13573_ net2496 net263 net396 vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10785_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[27\] net1041 vssd1
+ vssd1 vccd1 vccd1 _06782_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18100_ clknet_leaf_39_wb_clk_i _03423_ _01796_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_15312_ net1093 vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__inv_2
X_12524_ net1681 _03612_ net209 vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16292_ net1168 vssd1 vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18031_ clknet_leaf_97_wb_clk_i _03370_ _01727_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15243_ net1070 vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__inv_2
X_12455_ net1782 _03612_ net213 vssd1 vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__mux2_1
XANTENNA__12407__S net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11406_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[13\] _07328_
+ net1965 vssd1 vssd1 vccd1 vccd1 _07334_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15174_ net1247 vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__inv_2
X_12386_ net501 _07530_ _07796_ vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__a21o_2
XFILLER_0_23_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14125_ team_05_WB.instance_to_wrap.CPU_DAT_O\[12\] net507 _03858_ _03988_ vssd1
+ vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08964__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11337_ _07293_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.next_rows\[2\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_1_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_150_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_150_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_91_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13746__B _06521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14056_ _03901_ _03923_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11268_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[18\] _07125_
+ _07128_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[66\] vssd1 vssd1
+ vccd1 vccd1 _07229_ sky130_fd_sc_hd__a22o_1
X_13007_ _06423_ net2725 net460 vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__mux2_1
XANTENNA__13238__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08716__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10219_ _06102_ _06244_ vssd1 vssd1 vccd1 vccd1 _06245_ sky130_fd_sc_hd__or2_2
X_11199_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[54\] _07117_
+ _07120_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[38\] _07150_
+ vssd1 vssd1 vccd1 vccd1 _07164_ sky130_fd_sc_hd__a221o_1
XFILLER_0_158_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17815_ clknet_leaf_89_wb_clk_i _03158_ _01511_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[125\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09126__C1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13762__A net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17746_ clknet_leaf_95_wb_clk_i _03089_ _01442_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14958_ net1179 vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09141__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13909_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[26\]
+ net560 net576 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[26\]
+ net987 vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__a221o_1
XANTENNA__10287__B2 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17677_ clknet_leaf_102_wb_clk_i _03020_ _01373_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[115\]
+ sky130_fd_sc_hd__dfrtp_1
X_14889_ net1214 vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_46_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16628_ clknet_leaf_119_wb_clk_i _02258_ _00324_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09429__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16559_ clknet_leaf_133_wb_clk_i _02189_ _00255_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12984__A0 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09100_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[12\]
+ net694 net594 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[12\]
+ _05156_ vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__a221o_1
XFILLER_0_150_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09031_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[14\]
+ net823 _05087_ _05090_ vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__a211o_1
X_18229_ clknet_leaf_50_wb_clk_i net1457 _01924_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12544__C _03659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold301 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[91\] vssd1 vssd1
+ vccd1 vccd1 net1715 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold312 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[108\] vssd1 vssd1
+ vccd1 vccd1 net1726 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_27_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold323 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[28\] vssd1 vssd1
+ vccd1 vccd1 net1737 sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[63\] vssd1 vssd1
+ vccd1 vccd1 net1748 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08955__A2 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold345 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[114\] vssd1 vssd1
+ vccd1 vccd1 net1759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[9\] vssd1 vssd1
+ vccd1 vccd1 net1770 sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[46\] vssd1 vssd1
+ vccd1 vccd1 net1781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[65\] vssd1 vssd1
+ vccd1 vccd1 net1792 sky130_fd_sc_hd__dlygate4sd3_1
Xhold389 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[118\] vssd1 vssd1
+ vccd1 vccd1 net1803 sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ _05189_ _05825_ _05960_ _05937_ vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__a31o_1
XFILLER_0_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout803 net805 vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__buf_6
XFILLER_0_1_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout814 _04388_ vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__clkbuf_8
Xfanout825 _04384_ vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__buf_4
XANTENNA__11457__A net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13148__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08707__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout398_A _03731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout836 _04381_ vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__clkbuf_8
X_09864_ _04757_ _04799_ _05889_ _04756_ vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__o211a_1
Xfanout847 _04373_ vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__clkbuf_8
Xfanout858 net859 vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09572__D net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout869 net870 vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__buf_2
Xhold1001 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net2415 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1012 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net2426 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09380__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08815_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[18\]
+ net676 net625 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[18\]
+ _04883_ vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__a221o_1
Xhold1023 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net2437 sky130_fd_sc_hd__dlygate4sd3_1
X_09795_ _05823_ _05825_ vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__and2_1
XANTENNA__12987__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1034 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1045 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 net2459 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1056 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net2470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2481 sky130_fd_sc_hd__dlygate4sd3_1
X_08746_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[21\]
+ net717 _04813_ _04817_ vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__o22ai_4
Xhold1078 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[11\] vssd1
+ vssd1 vccd1 vccd1 net2492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1089 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2503 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout732_A _07030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08677_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[23\]
+ net843 net784 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout353_X net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11227__B1 _07127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout618_X net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_66_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13611__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10570_ _05237_ _06578_ _06051_ vssd1 vssd1 vccd1 vccd1 _06579_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09840__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09229_ net570 net534 _05260_ vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09747__D net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12240_ _03523_ _03526_ _03534_ _03520_ vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12171_ _07968_ _07972_ _07979_ _07971_ vssd1 vssd1 vccd1 vccd1 _07983_ sky130_fd_sc_hd__o22ai_2
XPHY_EDGE_ROW_2_Left_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10753__A2 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11122_ _07087_ _07088_ _07077_ vssd1 vssd1 vccd1 vccd1 _07089_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_82_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold890 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2304 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13058__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18211__Q team_05_WB.instance_to_wrap.total_design.core.instr_fetch vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15930_ net1289 vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__inv_2
X_11053_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[2\] net1044 net960
+ _07020_ vssd1 vssd1 vccd1 vccd1 _07021_ sky130_fd_sc_hd__o31a_1
XANTENNA__09108__Y _05165_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10004_ _06017_ _06032_ net372 vssd1 vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09371__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15861_ net1265 vssd1 vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__inv_2
XANTENNA__12897__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17600_ clknet_leaf_78_wb_clk_i _02971_ _01296_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_14812_ net1095 vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__inv_2
X_15792_ net1275 vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__inv_2
XANTENNA__09659__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17531_ clknet_leaf_80_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[2\]
+ _01227_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09123__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10269__B2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[26\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14743_ net1096 vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11955_ net343 _07761_ _07751_ net501 vssd1 vssd1 vccd1 vccd1 _07767_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_87_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08331__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17462_ clknet_leaf_59_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[30\]
+ _01158_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10906_ _06214_ _06768_ _06898_ _06900_ net568 vssd1 vssd1 vccd1 vccd1 _06901_ sky130_fd_sc_hd__a221o_1
X_14674_ net1238 vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11886_ _07689_ _07695_ _07697_ vssd1 vssd1 vccd1 vccd1 _07698_ sky130_fd_sc_hd__a21oi_2
X_16413_ clknet_leaf_108_wb_clk_i _02043_ _00109_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13625_ _04256_ net557 _03694_ vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__and3_4
X_17393_ clknet_leaf_65_wb_clk_i net1435 _01089_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10837_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[4\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06834_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13521__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15302__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16344_ clknet_leaf_27_wb_clk_i _01974_ _00040_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13556_ net1904 net323 net401 vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__mux2_1
X_10768_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[0\] net904 _04247_
+ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[0\] _06765_ vssd1 vssd1
+ vccd1 vccd1 _06766_ sky130_fd_sc_hd__a221o_1
XANTENNA__09831__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17497__Q team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10977__C1 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12507_ net1666 _03623_ net210 vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16275_ net1129 vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__inv_2
XANTENNA__10446__A net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13487_ net315 net2835 net411 vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__mux2_1
X_10699_ _06692_ _06693_ _06700_ net537 vssd1 vssd1 vccd1 vccd1 _06701_ sky130_fd_sc_hd__a31o_1
XFILLER_0_70_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18014_ clknet_leaf_82_wb_clk_i _03353_ _01710_ vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__dfrtp_1
XANTENNA__13915__C1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_46 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15226_ net1055 vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__inv_2
XFILLER_0_164_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12438_ _07847_ net919 vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_130_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08398__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08937__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15157_ net1061 vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12369_ net354 _03642_ _03626_ vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_50_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14108_ _04160_ _03950_ _04159_ vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__a21o_1
X_18374__1359 vssd1 vssd1 vccd1 vccd1 _18374__1359/HI net1359 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_39_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15088_ net1183 vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_39_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09673__C net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09347__C1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14039_ _03907_ _03908_ _03858_ vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__a21o_1
XANTENNA__11708__C team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[14\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire533_A _05575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09362__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08600_ net570 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[25\]
+ _04362_ vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__o21a_1
XANTENNA__12600__S _03680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13446__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09580_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[2\]
+ net940 net935 net926 vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__and4_1
XANTENNA__09114__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08531_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[26\]
+ net654 net641 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[26\]
+ _04607_ vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__a221o_1
X_17729_ clknet_leaf_98_wb_clk_i _03072_ _01425_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_100_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08462_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[28\]
+ net820 net765 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[28\]
+ _04540_ vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__a221o_1
XFILLER_0_174_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11209__B1 _07128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08393_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[29\]
+ net708 net658 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_102_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10680__B2 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13431__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09822__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_171_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1055_A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09567__D net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09014_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[14\]
+ net658 net635 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[14\]
+ _05064_ vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold120 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[7\]
+ vssd1 vssd1 vccd1 vccd1 net1534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[17\]
+ vssd1 vssd1 vccd1 vccd1 net1545 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold142 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[10\]
+ vssd1 vssd1 vccd1 vccd1 net1556 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1222_A net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold153 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[13\]
+ vssd1 vssd1 vccd1 vccd1 net1567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[8\]
+ vssd1 vssd1 vccd1 vccd1 net1578 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[10\]
+ vssd1 vssd1 vccd1 vccd1 net1589 sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[15\]
+ vssd1 vssd1 vccd1 vccd1 net1600 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09583__C net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout682_A _04301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold197 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[19\]
+ vssd1 vssd1 vccd1 vccd1 net1611 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout600 net601 vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__buf_4
Xfanout611 _04319_ vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout622 net624 vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__clkbuf_8
X_09916_ net517 _05731_ vssd1 vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout1010_X net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout633 _04313_ vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__buf_4
Xfanout644 net647 vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1108_X net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout655 _04308_ vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__buf_4
XFILLER_0_95_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09880__A _04573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout666 _04305_ vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__clkbuf_8
Xfanout677 net679 vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__clkbuf_8
X_09847_ _05871_ _05873_ _05875_ _05877_ vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__or4_1
Xfanout688 net690 vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout470_X net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout699 _04293_ vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout947_A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout568_X net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13606__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12510__S _03676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ _05508_ _05808_ _05506_ vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_126_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09105__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11634__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08729_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[21\]
+ net692 net645 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout735_X net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11740_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[9\] net997 vssd1
+ vssd1 vccd1 vccd1 _07552_ sky130_fd_sc_hd__nand2_2
XFILLER_0_138_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_189_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_37_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11671_ _06772_ _07485_ vssd1 vssd1 vccd1 vccd1 _07486_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout902_X net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13341__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12948__A0 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13410_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[16\]
+ net268 net416 vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10622_ net516 _06127_ _06129_ _06627_ vssd1 vssd1 vccd1 vccd1 _06628_ sky130_fd_sc_hd__a31oi_1
X_14390_ net1525 vssd1 vssd1 vccd1 vccd1 _02986_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_12_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09813__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09758__C net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13341_ net255 net2817 net424 vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10553_ net1018 _05187_ net551 _06562_ vssd1 vssd1 vccd1 vccd1 _06563_ sky130_fd_sc_hd__o31a_1
X_16060_ net1262 vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13272_ net229 net2206 net434 vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__mux2_1
X_10484_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[16\] net903 net965
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[16\] _06497_ vssd1
+ vssd1 vccd1 vccd1 _06498_ sky130_fd_sc_hd__a221o_1
XFILLER_0_161_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15011_ net1206 vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__inv_2
X_12223_ net547 _07751_ vssd1 vssd1 vccd1 vccd1 _03518_ sky130_fd_sc_hd__and2_2
XANTENNA__09041__A1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09774__B _05596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12154_ _07957_ _07965_ _07958_ vssd1 vssd1 vccd1 vccd1 _07966_ sky130_fd_sc_hd__o21a_1
XANTENNA__08154__A_N net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11105_ _07036_ _07070_ vssd1 vssd1 vccd1 vccd1 _07072_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_120_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16962_ clknet_leaf_5_wb_clk_i _02592_ _00658_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12085_ _07892_ _07896_ vssd1 vssd1 vccd1 vccd1 _07897_ sky130_fd_sc_hd__nor2_1
XANTENNA__09344__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15913_ net1270 vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__inv_2
X_11036_ _06832_ _06833_ _06849_ _07006_ vssd1 vssd1 vccd1 vccd1 _07007_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_34_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16893_ clknet_leaf_109_wb_clk_i _02523_ _00589_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13516__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15844_ net1299 vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__inv_2
XANTENNA__12420__S net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11439__B1 team_05_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15775_ net1293 vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12987_ _06655_ net2297 net466 vssd1 vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08304__B1 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17514_ clknet_leaf_73_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[17\]
+ _01210_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[17\]
+ sky130_fd_sc_hd__dfrtp_4
X_14726_ net1280 vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11938_ net501 _07527_ vssd1 vssd1 vccd1 vccd1 _07750_ sky130_fd_sc_hd__nor2_2
XFILLER_0_86_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17445_ clknet_leaf_60_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[13\]
+ _01141_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14657_ net1236 vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09949__B _05886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11869_ _07597_ _07680_ _07678_ vssd1 vssd1 vccd1 vccd1 _07681_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_60_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13251__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13608_ net2714 _06499_ net392 vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__mux2_1
X_17376_ clknet_leaf_64_wb_clk_i net1423 _01072_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14588_ net1083 vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09668__C net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16327_ net1119 vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13539_ net2349 net258 net400 vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__mux2_1
XANTENNA__09280__A1 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16258_ net1113 vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15209_ net1214 vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__inv_2
X_16189_ net1145 vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08791__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11438__C team_05_WB.instance_to_wrap.total_design.core.instr_fetch vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09701_ net512 _05731_ vssd1 vssd1 vccd1 vccd1 _05734_ sky130_fd_sc_hd__or2_1
XANTENNA__09335__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08543__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13426__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_74_Left_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09632_ net527 net523 vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_104_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09205__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[30\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09563_ _05599_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[2\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_172_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08514_ _04579_ _04587_ _04591_ net592 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[27\]
+ sky130_fd_sc_hd__o32a_4
XFILLER_0_148_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09494_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[4\]
+ net701 net645 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[4\]
+ _05532_ vssd1 vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08445_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[28\]
+ net674 net619 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[28\]
+ _04523_ vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout430_A net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_173_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16038__A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13161__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08376_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[30\]
+ net799 net734 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__a22o_1
XANTENNA__09578__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15877__A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_83_Left_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08074__A2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[24\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout316_X net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13355__A0 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11469__X _07380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout897_A net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12505__S _03673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1225_X net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout685_X net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08782__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout430 net431 vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__clkbuf_8
Xfanout441 _03716_ vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout452 net453 vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09326__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout463 _03711_ vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_92_Left_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout852_X net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout474 _03706_ vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__buf_6
XANTENNA__13336__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout485 _03703_ vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__buf_4
X_12910_ _06499_ net2644 net472 vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_6_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout496 net499 vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__buf_6
X_13890_ net1552 net981 _03781_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[16\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__10341__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12841_ net258 net2676 net481 vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ net1123 vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__inv_2
X_12772_ net254 net2493 net488 vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14511_ net1239 vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__inv_2
XANTENNA__10644__A1 _05577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11723_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[11\] net999 vssd1
+ vssd1 vccd1 vccd1 _07535_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15491_ net1171 vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18373__1358 vssd1 vssd1 vccd1 vccd1 _18373__1358/HI net1358 sky130_fd_sc_hd__conb_1
XFILLER_0_167_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13071__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17230_ clknet_leaf_177_wb_clk_i _02860_ _00926_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14442_ net1122 vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__inv_2
X_11654_ net8 net989 net916 net2410 vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__o22a_1
XFILLER_0_166_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12397__A1 _03666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17161_ clknet_leaf_21_wb_clk_i _02791_ _00857_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10605_ _06580_ _06611_ net517 vssd1 vssd1 vccd1 vccd1 _06612_ sky130_fd_sc_hd__mux2_1
X_14373_ _04144_ _04145_ vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__nand2_1
X_11585_ net2009 net1005 _07365_ net357 vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16112_ net1134 vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13324_ net2664 net310 net428 vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10536_ _06049_ _06211_ _06545_ net335 _06546_ vssd1 vssd1 vccd1 vccd1 _06547_ sky130_fd_sc_hd__o221ai_2
X_17092_ clknet_leaf_178_wb_clk_i _02722_ _00788_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_59 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16043_ net1250 vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__inv_2
X_13255_ net319 net2346 net438 vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12415__S net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10467_ _05015_ _05837_ vssd1 vssd1 vccd1 vccd1 _06481_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_122_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12206_ _07990_ _07993_ _07997_ _08013_ _08016_ vssd1 vssd1 vccd1 vccd1 _08018_ sky130_fd_sc_hd__o311ai_4
XFILLER_0_122_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_57_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_36_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13186_ net319 net2795 net442 vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__mux2_1
X_10398_ net334 _06240_ _06414_ _06415_ vssd1 vssd1 vccd1 vccd1 _06416_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_36_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11372__A2 _06756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08773__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12137_ _07948_ _07946_ vssd1 vssd1 vccd1 vccd1 _07949_ sky130_fd_sc_hd__and2b_1
XFILLER_0_20_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17994_ clknet_leaf_83_wb_clk_i _03333_ _01690_ vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09317__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13754__B _06369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12068_ _07868_ _07879_ vssd1 vssd1 vccd1 vccd1 _07880_ sky130_fd_sc_hd__nor2_1
X_16945_ clknet_leaf_168_wb_clk_i _02575_ _00641_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08525__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11555__A _07379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13246__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11019_ net1045 _06636_ _06992_ net959 vssd1 vssd1 vccd1 vccd1 _06993_ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10332__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16876_ clknet_leaf_0_wb_clk_i _02506_ _00572_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09670__D net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15827_ net1301 vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15758_ net1297 vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14709_ net1060 vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15689_ net1159 vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__inv_2
XANTENNA__09679__B net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08230_ net886 net861 net859 vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__and3_4
X_17428_ clknet_leaf_56_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[28\]
+ _01124_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08161_ _04229_ _04242_ vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__nand2_1
X_17359_ clknet_leaf_37_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[23\]
+ _01055_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14129__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08092_ net1025 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[15\]
+ net971 _04195_ vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload40 clknet_leaf_189_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload40/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_28_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload51 clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload51/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__11548__A_N _07407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload62 clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload62/Y sky130_fd_sc_hd__inv_16
Xclkload73 clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload73/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_77_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload84 clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload84/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_11_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload95 clknet_leaf_57_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload95/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__09556__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08994_ net571 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[15\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[15\] vssd1 vssd1 vccd1
+ vccd1 _05055_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout1018_A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09308__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13156__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout478_A net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10323__B1 _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09580__D net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09615_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[2\]
+ net880 net870 net866 vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__and4_1
XFILLER_0_92_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout645_A net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09546_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[3\]
+ net687 net656 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[3\]
+ _05580_ vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10626__A1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09477_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[4\]
+ net834 net816 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[4\]
+ _05516_ vssd1 vssd1 vccd1 vccd1 _05517_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout812_A net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09492__A1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout433_X net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1175_X net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08428_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[29\]
+ net755 net738 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[29\]
+ _04507_ vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__a221o_1
XFILLER_0_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12379__A1 _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload1 clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload1/X sky130_fd_sc_hd__clkbuf_8
X_08359_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[30\]
+ net688 net657 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[30\]
+ _04439_ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout600_X net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15400__A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11370_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[1\] _07308_ _06769_
+ vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__mux2_1
XANTENNA__08452__C1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10321_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[24\] _06099_ vssd1
+ vssd1 vccd1 vccd1 _06343_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10544__A net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09755__D net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09547__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13040_ net252 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[20\]
+ net456 vssd1 vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__mux2_1
X_10252_ net894 _06275_ _06274_ net555 vssd1 vssd1 vccd1 vccd1 _06276_ sky130_fd_sc_hd__a211o_1
XANTENNA__08755__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10183_ _06208_ _06209_ net529 vssd1 vssd1 vccd1 vccd1 _06210_ sky130_fd_sc_hd__mux2_1
Xfanout1203 net1206 vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__buf_4
Xfanout1214 net1215 vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__buf_4
Xfanout1225 net1241 vssd1 vssd1 vccd1 vccd1 net1225 sky130_fd_sc_hd__buf_4
Xfanout1236 net1237 vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__buf_4
XANTENNA_input39_A wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08301__X _04383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14991_ net1282 vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__inv_2
Xfanout1247 net1252 vssd1 vssd1 vccd1 vccd1 net1247 sky130_fd_sc_hd__buf_4
Xfanout1258 net1261 vssd1 vssd1 vccd1 vccd1 net1258 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_31_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout260 net262 vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__buf_2
Xfanout1269 net1270 vssd1 vssd1 vccd1 vccd1 net1269 sky130_fd_sc_hd__buf_4
Xfanout271 net272 vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_31_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08507__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13066__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout282 net285 vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__buf_2
X_13942_ _03811_ _03815_ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__or2_1
X_16730_ clknet_leaf_31_wb_clk_i _02360_ _00426_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout293 _06588_ vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16661_ clknet_leaf_24_wb_clk_i _02291_ _00357_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13873_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[8\]
+ net559 net575 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[8\]
+ net986 vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_175_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_175_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15612_ net1150 vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18400_ net1372 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__buf_2
X_12824_ net309 net2590 net485 vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__mux2_1
X_16592_ clknet_leaf_167_wb_clk_i _02222_ _00288_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_104_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_104_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08684__A net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18331_ net1320 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
X_15543_ net1139 vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__inv_2
X_12755_ net329 net2530 net494 vssd1 vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11706_ net550 _07515_ vssd1 vssd1 vccd1 vccd1 _07518_ sky130_fd_sc_hd__nand2_2
X_18262_ clknet_leaf_37_wb_clk_i _03491_ _01957_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[16\]
+ sky130_fd_sc_hd__dfrtp_4
X_15474_ net1173 vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__inv_2
X_12686_ net2948 net339 vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__and2_1
XANTENNA__08971__X _05034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14425_ net1057 vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17213_ clknet_leaf_108_wb_clk_i _02843_ _00909_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11637_ team_05_WB.instance_to_wrap.BUSY_O net991 team_05_WB.instance_to_wrap.wishbone.prev_BUSY_O
+ vssd1 vssd1 vccd1 vccd1 _07484_ sky130_fd_sc_hd__or3b_1
X_18193_ clknet_leaf_34_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[14\]
+ _01888_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17144_ clknet_leaf_32_wb_clk_i _02774_ _00840_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14356_ _04098_ _04104_ _04103_ vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__o21ba_1
X_11568_ net920 _07354_ _07422_ net1007 net1582 vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__a32o_1
XANTENNA__13749__B _06464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13307_ net2479 net252 net428 vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__mux2_1
Xhold708 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 net2122 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11593__A2 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10519_ _06049_ _06141_ _06378_ _06503_ vssd1 vssd1 vccd1 vccd1 _06531_ sky130_fd_sc_hd__o22a_1
Xhold719 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2133 sky130_fd_sc_hd__dlygate4sd3_1
X_17075_ clknet_leaf_166_wb_clk_i _02705_ _00771_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14287_ _06350_ _04060_ _06918_ _06320_ vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_126_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11499_ _07404_ _07405_ _07407_ _07409_ _07402_ vssd1 vssd1 vccd1 vccd1 _07410_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_0_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_139_Left_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16026_ net1284 vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__inv_2
X_13238_ net232 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[23\]
+ net439 vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13169_ net230 net2609 net443 vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17977_ clknet_leaf_74_wb_clk_i _03316_ _01673_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__dfrtp_1
Xhold1408 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2822 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14295__A1 _04613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1419 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2833 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14295__B2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[25\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16928_ clknet_leaf_133_wb_clk_i _02558_ _00624_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09171__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16859_ clknet_leaf_191_wb_clk_i _02489_ _00555_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_140_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_148_Left_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09400_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[18\] net965
+ _04269_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[26\] _05444_
+ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[6\]
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10608__A1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09331_ _05376_ _05377_ vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__nor2_4
XFILLER_0_88_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09262_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[9\]
+ net772 net758 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08213_ _04232_ net962 _04271_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[17\]
+ _04153_ vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__o311a_2
XTAP_TAPCELL_ROW_138_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09193_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[10\]
+ net664 net629 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08144_ _04213_ _04224_ vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09777__A2 _05807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_157_Left_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08985__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload140 clknet_leaf_150_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload140/X sky130_fd_sc_hd__clkbuf_4
X_08075_ net1025 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__and2b_1
Xclkload151 clknet_leaf_136_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload151/Y sky130_fd_sc_hd__clkinv_4
XANTENNA_fanout1135_A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload162 clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload162/Y sky130_fd_sc_hd__inv_6
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09575__D net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload173 clknet_leaf_103_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload173/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_168_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload184 clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload184/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_144_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09529__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12533__A1 _03605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08737__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout595_A net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08201__A2 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18372__1357 vssd1 vssd1 vccd1 vccd1 _18372__1357/HI net1357 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_164_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold13 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[9\]
+ vssd1 vssd1 vccd1 vccd1 net1427 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[24\]
+ vssd1 vssd1 vccd1 vccd1 net1438 sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[15\]
+ net849 net752 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[15\]
+ _05038_ vssd1 vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__a221o_1
Xhold35 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[0\]
+ vssd1 vssd1 vccd1 vccd1 net1449 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout762_A net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout383_X net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold46 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[17\]
+ vssd1 vssd1 vccd1 vccd1 net1460 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold57 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[23\]
+ vssd1 vssd1 vccd1 vccd1 net1471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[28\]
+ vssd1 vssd1 vccd1 vccd1 net1482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[3\]
+ vssd1 vssd1 vccd1 vccd1 net1493 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09162__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_166_Left_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12578__X _03681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout648_X net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13614__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11923__A team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10870_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[16\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[16\]
+ _06866_ vssd1 vssd1 vccd1 vccd1 _06867_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09529_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[3\]
+ net774 net771 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[3\]
+ _05559_ vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout815_X net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12540_ net1883 _03641_ net209 vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1062 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10973__S net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12471_ net1792 _03641_ net213 vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14210_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[9\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[10\]
+ _04006_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[11\] vssd1
+ vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__a31o_1
XFILLER_0_151_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11422_ _04165_ _07321_ vssd1 vssd1 vccd1 vccd1 _07340_ sky130_fd_sc_hd__and2_1
X_15190_ net1091 vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__inv_2
XANTENNA__09768__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14141_ net2974 net506 net912 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[24\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__08976__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11353_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[4\] net508 _07296_
+ team_05_WB.instance_to_wrap.total_design.data_from_keypad\[0\] vssd1 vssd1 vccd1
+ vccd1 _03387_ sky130_fd_sc_hd__a22o_1
XANTENNA__10274__A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08440__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10304_ net525 _06223_ vssd1 vssd1 vccd1 vccd1 _06326_ sky130_fd_sc_hd__nand2_1
X_14072_ _03914_ _03918_ _03938_ _03939_ vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11284_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[50\] _07110_
+ _07230_ _07244_ vssd1 vssd1 vccd1 vccd1 _07245_ sky130_fd_sc_hd__a211o_1
XFILLER_0_104_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11327__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12524__A1 _03612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08728__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17900_ clknet_leaf_88_wb_clk_i _03243_ _01596_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13023_ net329 net2484 net462 vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__mux2_1
X_10235_ _06195_ _06259_ net521 vssd1 vssd1 vccd1 vccd1 _06260_ sky130_fd_sc_hd__mux2_1
Xfanout1000 _07470_ vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__buf_2
Xfanout1011 net1012 vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__clkbuf_4
X_17831_ clknet_leaf_87_wb_clk_i _03174_ _01527_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[77\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1022 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[6\] vssd1
+ vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__clkbuf_4
Xfanout1033 net1035 vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__clkbuf_4
X_10166_ net1020 _04512_ _04514_ net552 vssd1 vssd1 vccd1 vccd1 _06193_ sky130_fd_sc_hd__a211o_1
Xfanout1044 net1047 vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__buf_2
Xfanout1055 net1056 vssd1 vssd1 vccd1 vccd1 net1055 sky130_fd_sc_hd__buf_4
Xfanout1066 net1067 vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__buf_4
X_17762_ clknet_leaf_98_wb_clk_i _03105_ _01458_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1077 net1078 vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__buf_4
Xfanout1088 net1094 vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__buf_2
X_14974_ net1066 vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__inv_2
X_10097_ _06117_ _06124_ net526 vssd1 vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__mux2_2
Xfanout1099 net1100 vssd1 vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__buf_4
X_16713_ clknet_leaf_21_wb_clk_i _02343_ _00409_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13925_ net910 _03800_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[0\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17693_ clknet_leaf_92_wb_clk_i _03036_ _01389_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[67\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13524__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload4_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13856_ team_05_WB.instance_to_wrap.total_design.core.data_mem.state\[2\] _04177_
+ net726 team_05_WB.instance_to_wrap.total_design.core.data_mem.state\[0\] vssd1 vssd1
+ vccd1 vccd1 _03764_ sky130_fd_sc_hd__and4b_1
X_16644_ clknet_leaf_183_wb_clk_i _02274_ _00340_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12807_ net252 net2956 net484 vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13787_ _04171_ team_05_WB.instance_to_wrap.total_design.core.data_mem.state\[2\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.state\[1\] net726 vssd1 vssd1
+ vccd1 vccd1 _03760_ sky130_fd_sc_hd__or4_1
XANTENNA__12000__Y _07812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16575_ clknet_leaf_153_wb_clk_i _02205_ _00271_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08259__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10999_ net963 _06557_ _06976_ vssd1 vssd1 vccd1 vccd1 _06977_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18314_ net1406 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
X_15526_ net1158 vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__inv_2
X_12738_ net248 net2546 net494 vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15457_ net1156 vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__inv_2
X_18245_ clknet_leaf_52_wb_clk_i net1031 _01940_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.disable_pc_reg
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_44_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10736__X _06736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12669_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[20\]
+ net339 vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14408_ net1532 vssd1 vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11015__A1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09759__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_160_Right_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18176_ clknet_leaf_51_wb_clk_i net1614 _01871_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_72_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15388_ net1095 vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_96_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09676__C net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08206__X _04289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08967__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_64_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17127_ clknet_leaf_203_wb_clk_i _02757_ _00823_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_14339_ _05123_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[13\]
+ _05165_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__a22o_1
Xhold505 net92 vssd1 vssd1 vccd1 vccd1 net1919 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold516 net137 vssd1 vssd1 vccd1 vccd1 net1930 sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net1941 sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1952 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17058_ clknet_leaf_8_wb_clk_i _02688_ _00754_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold549 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1963 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11318__A2 _07091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08719__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08900_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[17\] vssd1
+ vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__inv_2
X_16009_ net1112 vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__inv_2
XANTENNA__12603__S _03681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09880_ _04573_ _04592_ vssd1 vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_111_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09392__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08831_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[18\]
+ net715 _04896_ _04899_ vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_100_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1205 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1216 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2630 sky130_fd_sc_hd__dlygate4sd3_1
X_08762_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[21\]
+ net830 net791 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[21\]
+ _04833_ vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__a221o_1
Xhold1227 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2641 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1238 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2652 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1249 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2663 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09144__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08498__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08693_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[22\]
+ net681 net631 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__a22o_1
XANTENNA__13434__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1085_A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09314_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[8\]
+ net828 net824 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_56_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_48_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09245_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[9\]
+ net701 net608 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout510_A net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08670__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1252_A net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout608_A _04320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09176_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[11\]
+ net782 net756 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[11\]
+ _05217_ vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08958__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08127_ net152 net151 vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__nand2_1
XANTENNA__08422__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08058_ _04171_ team_05_WB.instance_to_wrap.total_design.core.data_mem.state\[2\]
+ _04177_ vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__and3_1
XFILLER_0_141_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11309__A2 _07109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12506__A1 _03641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout598_X net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13609__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12513__S net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10517__B1 _06160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10020_ _05531_ _06002_ vssd1 vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__or2_4
XANTENNA__09383__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11637__B net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11190__B1 _07100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout765_X net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09135__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_95_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10968__S net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11971_ _07726_ _07743_ _07728_ vssd1 vssd1 vccd1 vccd1 _07783_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout932_X net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08489__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13710_ net901 _06591_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[10\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__13344__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10922_ net1044 _06291_ vssd1 vssd1 vccd1 vccd1 _06914_ sky130_fd_sc_hd__nor2_1
X_14690_ net1226 vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__inv_2
X_13641_ net2284 net268 net388 vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__mux2_1
X_10853_ _06833_ _06849_ _06832_ vssd1 vssd1 vccd1 vccd1 _06850_ sky130_fd_sc_hd__a21bo_1
X_16360_ clknet_leaf_196_wb_clk_i _01990_ _00056_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13572_ net2315 net255 net396 vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10784_ _06779_ _06780_ vssd1 vssd1 vccd1 vccd1 _06781_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15311_ net1233 vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__inv_2
X_12523_ net1881 _03614_ net209 vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16291_ net1164 vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_23_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18030_ clknet_leaf_97_wb_clk_i _03369_ _01726_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_15242_ net1122 vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__inv_2
X_12454_ net1786 _03614_ net213 vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11405_ _07330_ _07333_ vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15173_ net1194 vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__inv_2
X_12385_ net1766 _07812_ _07852_ vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_202_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08413__A2 _04417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14124_ _03985_ _03986_ vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__xnor2_1
X_11336_ net152 net151 net154 net153 vssd1 vssd1 vccd1 vccd1 _07293_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_91_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13519__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14055_ _03901_ _03923_ vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__or2_1
X_11267_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[42\] _07091_
+ _07109_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[74\] vssd1 vssd1
+ vccd1 vccd1 _07228_ sky130_fd_sc_hd__a22o_1
XANTENNA__12423__S _03667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09374__B1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13006_ net246 net2931 net462 vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__mux2_1
X_10218_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[27\] _06101_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[28\]
+ vssd1 vssd1 vccd1 vccd1 _06244_ sky130_fd_sc_hd__a21oi_1
X_11198_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[126\] _07099_
+ _07109_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[78\] _07162_
+ vssd1 vssd1 vccd1 vccd1 _07163_ sky130_fd_sc_hd__a221o_1
XANTENNA__11181__B1 _07106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_190_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_190_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_118_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17814_ clknet_leaf_76_wb_clk_i _03157_ _01510_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[124\]
+ sky130_fd_sc_hd__dfrtp_1
X_10149_ net524 _06170_ _06176_ net333 vssd1 vssd1 vccd1 vccd1 _06177_ sky130_fd_sc_hd__a211o_1
XFILLER_0_89_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13762__B _06108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17745_ clknet_leaf_98_wb_clk_i _03088_ _01441_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[55\]
+ sky130_fd_sc_hd__dfrtp_1
X_14957_ net1081 vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13254__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13908_ net1546 net983 _03790_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[25\]
+ sky130_fd_sc_hd__o21a_1
X_17676_ clknet_leaf_77_wb_clk_i _03019_ _01372_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[114\]
+ sky130_fd_sc_hd__dfrtp_1
X_14888_ net1216 vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16627_ clknet_leaf_166_wb_clk_i _02257_ _00323_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13839_ net1460 net579 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[17\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16558_ clknet_leaf_177_wb_clk_i _02188_ _00254_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18371__1356 vssd1 vssd1 vccd1 vccd1 _18371__1356/HI net1356 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_21_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15509_ net1172 vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_21_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12394__A _07864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08652__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16489_ clknet_leaf_22_wb_clk_i _02119_ _00185_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11502__S net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09030_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[14\]
+ net842 _05088_ _05089_ vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__a211o_1
X_18228_ clknet_leaf_57_wb_clk_i net1605 _01923_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18159_ clknet_leaf_167_wb_clk_i _03462_ _01855_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold302 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1716 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold313 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[66\] vssd1 vssd1
+ vccd1 vccd1 net1727 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold324 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[56\] vssd1 vssd1
+ vccd1 vccd1 net1738 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10340__A1_N _05924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold335 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[124\] vssd1 vssd1
+ vccd1 vccd1 net1749 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold346 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[109\] vssd1 vssd1
+ vccd1 vccd1 net1760 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold357 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[52\] vssd1 vssd1
+ vccd1 vccd1 net1771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold368 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[81\] vssd1 vssd1
+ vccd1 vccd1 net1782 sky130_fd_sc_hd__dlygate4sd3_1
X_09932_ _05825_ _05960_ vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__nand2_1
XANTENNA__13429__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold379 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[50\] vssd1 vssd1
+ vccd1 vccd1 net1793 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout804 net805 vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__buf_2
XANTENNA__09365__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout815 _04388_ vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09208__A _05260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout826 _04383_ vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__buf_6
XFILLER_0_110_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09863_ _04756_ _04798_ vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__and2_1
Xfanout837 net840 vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__buf_6
Xfanout848 _04373_ vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__buf_4
XANTENNA__11172__B1 _07121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout293_A _06588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout859 _04298_ vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__clkbuf_4
Xhold1002 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2416 sky130_fd_sc_hd__dlygate4sd3_1
X_08814_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[18\]
+ net652 net621 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__a22o_1
Xhold1013 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2427 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1000_A _07470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09794_ _05208_ _05236_ vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__or2_1
Xhold1024 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net2438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1035 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net2449 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09117__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1046 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2460 sky130_fd_sc_hd__dlygate4sd3_1
X_08745_ _04802_ _04805_ _04815_ _04816_ vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__or4_1
Xhold1057 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net2471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1068 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2482 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout460_A _03711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1079 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 net2493 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout558_A net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13164__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08676_ _04743_ _04745_ _04747_ _04749_ vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_159_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_179_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout725_A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout346_X net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08891__A2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10986__B1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09228_ net534 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[10\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_1_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09159_ _04233_ net958 net921 _04147_ vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__a31o_1
XFILLER_0_82_1010 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12170_ _07936_ _07940_ _07979_ _07980_ _07931_ vssd1 vssd1 vccd1 vccd1 _07982_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_32_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13847__B net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout882_X net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11121_ _07063_ _07065_ vssd1 vssd1 vccd1 vccd1 _07088_ sky130_fd_sc_hd__nand2_1
XANTENNA__13339__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold880 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[0\]
+ vssd1 vssd1 vccd1 vccd1 net2305 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09356__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11052_ _06844_ _06899_ _07019_ vssd1 vssd1 vccd1 vccd1 _07020_ sky130_fd_sc_hd__or3b_1
X_10003_ _06024_ _06031_ net530 vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__mux2_1
X_15860_ net1299 vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__inv_2
XANTENNA__14311__X _04084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input21_A DAT_I[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14811_ net1078 vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__inv_2
X_15791_ net1294 vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13074__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17530_ clknet_leaf_66_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[1\]
+ _01226_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10269__A2 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11954_ net343 _07761_ vssd1 vssd1 vccd1 vccd1 _07766_ sky130_fd_sc_hd__nand2_1
X_14742_ net1084 vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10905_ _06884_ _06897_ vssd1 vssd1 vccd1 vccd1 _06900_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_28_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17461_ clknet_leaf_60_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[29\]
+ _01157_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_14673_ net1189 vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11885_ _07655_ _07696_ _07662_ vssd1 vssd1 vccd1 vccd1 _07697_ sky130_fd_sc_hd__o21a_1
XFILLER_0_15_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output108_A net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08882__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_103_Left_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12415__A0 _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16412_ clknet_leaf_157_wb_clk_i _02042_ _00108_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13624_ net2343 net306 net393 vssd1 vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__mux2_1
X_10836_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[5\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06833_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17392_ clknet_leaf_61_wb_clk_i net1438 _01088_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16343_ net1147 vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__inv_2
X_13555_ net2185 net311 net400 vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12418__S _03668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10767_ net536 _06764_ vssd1 vssd1 vccd1 vccd1 _06765_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_41_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12506_ net1836 _03641_ net211 vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__mux2_1
X_16274_ net1115 vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__inv_2
X_13486_ net317 net2475 net409 vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__mux2_1
X_10698_ net334 _06225_ net332 _06561_ _06699_ vssd1 vssd1 vccd1 vccd1 _06700_ sky130_fd_sc_hd__o221a_1
XFILLER_0_54_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10446__B _06461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18013_ clknet_leaf_82_wb_clk_i _03352_ _01709_ vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_164_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15225_ net1051 vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__inv_2
X_12437_ _03623_ net1789 net215 vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13391__A1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15156_ net1075 vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13757__B _06918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12368_ net1661 _03661_ net216 vssd1 vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10154__A2_N _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12661__B net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14107_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[15\] net978 _04159_
+ _04160_ vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__o211ai_2
XPHY_EDGE_ROW_112_Left_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13249__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11319_ _07272_ _07275_ _07276_ _07277_ vssd1 vssd1 vccd1 vccd1 _07278_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15087_ net1282 vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__inv_2
X_12299_ _03592_ _03593_ _03575_ vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_39_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09673__D net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08203__Y _04286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14038_ _03877_ _03879_ _03906_ vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__nand3_1
XANTENNA__14340__B1 _05256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13694__A2 _07349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15989_ net1128 vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08530_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[26\]
+ net685 net650 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__a22o_1
X_17728_ clknet_leaf_93_wb_clk_i _03071_ _01424_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_65_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_121_Left_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08461_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[28\]
+ net811 net769 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17659_ clknet_leaf_76_wb_clk_i _03002_ _01355_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[97\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08873__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12406__A0 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08392_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[29\]
+ net687 net605 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_102_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10968__A0 _06445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08625__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_171_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09013_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[14\]
+ net596 _05073_ net721 vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_171_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout306_A net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold110 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[4\] vssd1 vssd1
+ vccd1 vccd1 net1524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.state\[1\] vssd1 vssd1
+ vccd1 vccd1 net1535 sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[25\]
+ vssd1 vssd1 vccd1 vccd1 net1546 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09050__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold143 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[12\]
+ vssd1 vssd1 vccd1 vccd1 net1557 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[24\]
+ vssd1 vssd1 vccd1 vccd1 net1568 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13159__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold165 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[13\]
+ vssd1 vssd1 vccd1 vccd1 net1579 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[18\]
+ vssd1 vssd1 vccd1 vccd1 net1590 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1215_A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09583__D net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold187 net121 vssd1 vssd1 vccd1 vccd1 net1601 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09338__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout601 _04322_ vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__clkbuf_8
Xfanout612 _04319_ vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__clkbuf_8
Xhold198 net110 vssd1 vssd1 vccd1 vccd1 net1612 sky130_fd_sc_hd__dlygate4sd3_1
X_09915_ net366 _05801_ vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__or2_1
Xfanout623 net624 vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__buf_4
XANTENNA__12998__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout634 net635 vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__clkbuf_8
Xfanout645 net647 vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__clkbuf_8
Xfanout656 net659 vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__clkbuf_8
X_09846_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[20\]
+ net845 _05876_ net853 vssd1 vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__a211o_1
Xfanout667 _04305_ vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12893__A0 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1003_X net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout678 net679 vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__buf_4
Xfanout689 net690 vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__buf_4
X_09777_ _05552_ _05807_ _05551_ vssd1 vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_126_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout463_X net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout842_A net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08728_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[21\]
+ net673 net615 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__a22o_1
XANTENNA__08849__C1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout630_X net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08659_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[23\]
+ net706 net657 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[23\]
+ _04721_ vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_1_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08864__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13622__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11670_ net1050 team_05_WB.instance_to_wrap.total_design.core.instr_fetch vssd1 vssd1
+ vccd1 vccd1 _07485_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10621_ net513 _06126_ _06137_ vssd1 vssd1 vccd1 vccd1 _06627_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09758__D net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09895__X _05924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13340_ net252 net2947 net424 vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10552_ _05186_ _06051_ net511 _05189_ vssd1 vssd1 vccd1 vccd1 _06562_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__11620__B2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[10\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13271_ net233 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[23\]
+ net435 vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__mux2_1
X_10483_ net896 _06496_ vssd1 vssd1 vccd1 vccd1 _06497_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_129_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_129_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15010_ net1219 vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__inv_2
X_12222_ _07774_ net355 vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input69_A wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09041__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[14\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13069__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12153_ _07950_ _07953_ vssd1 vssd1 vccd1 vccd1 _07965_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11104_ _07036_ _07070_ vssd1 vssd1 vccd1 vccd1 _07071_ sky130_fd_sc_hd__and2b_1
X_12084_ _07884_ _07888_ _07890_ vssd1 vssd1 vccd1 vccd1 _07896_ sky130_fd_sc_hd__and3_1
X_16961_ clknet_leaf_150_wb_clk_i _02591_ _00657_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11528__D _07438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11035_ net1046 _07005_ vssd1 vssd1 vccd1 vccd1 _07006_ sky130_fd_sc_hd__nand2_1
X_15912_ net1265 vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__inv_2
X_18370__1355 vssd1 vssd1 vccd1 vccd1 _18370__1355/HI net1355 sky130_fd_sc_hd__conb_1
XANTENNA__12701__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16892_ clknet_leaf_159_wb_clk_i _02522_ _00588_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15843_ net1304 vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11439__A1 _07349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12636__A0 _03605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15774_ net1273 vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__inv_2
X_12986_ net294 net2828 net467 vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__mux2_1
XANTENNA__09501__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17513_ clknet_leaf_113_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[16\]
+ _01209_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_14725_ net1185 vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__inv_2
X_11937_ _07748_ vssd1 vssd1 vccd1 vccd1 _07749_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13532__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17444_ clknet_leaf_60_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[12\]
+ _01140_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10662__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11868_ _07648_ _07678_ _07641_ vssd1 vssd1 vccd1 vccd1 _07680_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14656_ net1200 vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10819_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[12\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06816_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13607_ net2464 net262 net393 vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17375_ clknet_leaf_81_wb_clk_i net1432 _01071_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08607__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14587_ net1098 vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__inv_2
X_11799_ _07589_ _07596_ vssd1 vssd1 vccd1 vccd1 _07611_ sky130_fd_sc_hd__xor2_2
XANTENNA__09668__D net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16326_ net1123 vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13538_ net2253 net254 net400 vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09280__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16257_ net1133 vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__inv_2
X_13469_ net233 net2839 net411 vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__mux2_1
XANTENNA__10744__X _06743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15208_ net1217 vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__inv_2
X_16188_ net1145 vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09684__C net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09032__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15139_ net1200 vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__inv_2
XANTENNA__09981__A net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17971__Q net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09700_ net512 _05731_ vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_147_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09631_ _05662_ _05664_ _05665_ _05635_ vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__o31ai_2
XANTENNA__12627__A0 _03612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09562_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[14\] net966
+ _04267_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[22\] _05598_
+ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__a221oi_1
XTAP_TAPCELL_ROW_104_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09099__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08513_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[27\]
+ net838 _04588_ _04590_ net855 vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_19_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09493_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[4\]
+ net677 net669 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08846__A2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout256_A _06442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13442__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08444_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[28\]
+ net714 net709 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_173_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08375_ _04449_ _04451_ _04453_ _04455_ vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout1165_A net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09578__D net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09271__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout211_X net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09023__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout792_A net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14304__B1 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout580_X net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout420 net423 vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__buf_6
XANTENNA_fanout678_X net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout431 _03723_ vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__buf_6
XANTENNA__11485__X _07396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13617__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout442 _03716_ vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__buf_6
XANTENNA__12521__S net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout453 _03713_ vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__buf_4
Xfanout464 _03710_ vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__buf_6
XANTENNA__14302__A _04533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout475 _03706_ vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__buf_4
Xfanout486 _03703_ vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_6_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout497 net499 vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__buf_6
X_09829_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[20\]
+ net715 _05856_ _05859_ vssd1 vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__o22ai_4
XANTENNA_fanout845_X net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12840_ net252 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[20\]
+ net480 vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08298__B1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[21\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12771_ net246 net2780 net490 vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08837__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13352__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11722_ _07479_ _07530_ vssd1 vssd1 vccd1 vccd1 _07534_ sky130_fd_sc_hd__nor2_1
X_14510_ net1188 vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__inv_2
X_15490_ net1167 vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_81_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11841__B2 _07623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1082 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09131__A _05165_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13043__A0 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14441_ net1214 vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__inv_2
X_11653_ net9 net989 net916 net2298 vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__o22a_1
X_10604_ _06019_ _06021_ vssd1 vssd1 vccd1 vccd1 _06611_ sky130_fd_sc_hd__nand2_1
X_14372_ net511 _06061_ _04142_ vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__mux2_1
X_17160_ clknet_leaf_204_wb_clk_i _02790_ _00856_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11584_ net2053 net1005 _07363_ net357 vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09262__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16111_ net1134 vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13323_ net2034 net330 net429 vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10535_ net1018 _05145_ _05830_ net551 vssd1 vssd1 vccd1 vccd1 _06546_ sky130_fd_sc_hd__a211o_1
XFILLER_0_88_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17091_ clknet_leaf_198_wb_clk_i _02721_ _00787_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08470__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16042_ net1287 vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__inv_2
X_13254_ net302 net2554 net438 vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10466_ net2543 net262 net542 vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__mux2_1
XANTENNA__09014__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12205_ _07990_ _07993_ _07997_ _08013_ vssd1 vssd1 vccd1 vccd1 _08017_ sky130_fd_sc_hd__o31a_1
XANTENNA__08758__D1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13185_ net303 net2038 net442 vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10397_ net337 _06228_ _06355_ _06225_ vssd1 vssd1 vccd1 vccd1 _06415_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_36_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_6_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_36_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12136_ _07881_ _07942_ vssd1 vssd1 vccd1 vccd1 _07948_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17993_ clknet_leaf_82_wb_clk_i _03332_ _01689_ vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__dfrtp_1
XANTENNA__13527__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12431__S net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12067_ _07865_ _07876_ _07874_ vssd1 vssd1 vccd1 vccd1 _07879_ sky130_fd_sc_hd__a21oi_1
X_16944_ clknet_leaf_138_wb_clk_i _02574_ _00640_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15308__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_97_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_53_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11018_ _06827_ _06852_ _06853_ _06991_ _04170_ vssd1 vssd1 vccd1 vccd1 _06992_ sky130_fd_sc_hd__a311o_1
XANTENNA__11555__B _07465_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_26_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16875_ clknet_leaf_188_wb_clk_i _02505_ _00571_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12609__A0 _03641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15826_ net1290 vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_142_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15757_ net1290 vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__inv_2
XANTENNA__08828__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12969_ net238 net2709 net466 vssd1 vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14708_ net1067 vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15688_ net1171 vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__inv_2
XANTENNA__09679__C net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08209__X _04292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17427_ clknet_leaf_66_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[27\]
+ _01123_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_145_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14639_ net1239 vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08160_ _04229_ _04242_ vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__and2_1
X_17358_ clknet_leaf_33_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[22\]
+ _01054_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10399__A1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11596__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16309_ net1160 vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08461__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08091_ net1025 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__and2b_1
XANTENNA__12606__S _03680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17289_ clknet_leaf_25_wb_clk_i _02919_ _00985_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11510__S net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire381_X net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload30 clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload30/Y sky130_fd_sc_hd__clkinv_8
Xclkload41 clknet_leaf_190_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload41/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_70_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10193__Y _06219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload52 clknet_leaf_174_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload52/Y sky130_fd_sc_hd__inv_6
XANTENNA__09005__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload63 clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload63/Y sky130_fd_sc_hd__inv_12
Xclkload74 clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload74/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_77_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload85 clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload85/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_101_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload96 clknet_leaf_58_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload96/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_149_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08993_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[15\]
+ net590 _05045_ _05054_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[15\]
+ sky130_fd_sc_hd__o22a_4
XFILLER_0_142_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13437__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10323__A1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[24\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10323__B2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[24\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09614_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[2\]
+ net877 net864 net862 vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__and4_1
X_09545_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[3\]
+ net664 net602 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[3\]
+ _05581_ vssd1 vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout540_A net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08819__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13172__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout259_X net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout638_A _04312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_174_Right_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09476_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[4\]
+ net753 net734 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__a22o_1
XANTENNA__10368__Y _06387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09492__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13025__A0 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08427_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[29\]
+ _04366_ net822 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[29\]
+ net854 vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__a221o_1
XFILLER_0_148_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14792__A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout426_X net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09886__A _04533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08358_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[30\]
+ net701 net634 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload2 clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload2/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__09244__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12516__S net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10384__X _06403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08289_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[23\] team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10320_ net537 _06341_ vssd1 vssd1 vccd1 vccd1 _06342_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13879__A2 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10544__B _06554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout795_X net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10251_ _04637_ _05991_ vssd1 vssd1 vccd1 vccd1 _06275_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09892__Y _05921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08789__X team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[19\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13855__B net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10182_ _06020_ _06030_ net519 vssd1 vssd1 vccd1 vccd1 _06209_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout962_X net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1204 net1206 vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__buf_4
Xfanout1215 net1241 vssd1 vssd1 vccd1 vccd1 net1215 sky130_fd_sc_hd__buf_4
XANTENNA__13347__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1226 net1234 vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__buf_4
Xfanout1237 net1241 vssd1 vssd1 vccd1 vccd1 net1237 sky130_fd_sc_hd__clkbuf_2
X_14990_ net1190 vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__inv_2
Xfanout1248 net1252 vssd1 vssd1 vccd1 vccd1 net1248 sky130_fd_sc_hd__buf_4
Xfanout1259 net1261 vssd1 vssd1 vccd1 vccd1 net1259 sky130_fd_sc_hd__buf_4
XANTENNA__09704__B1 _05212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout261 net262 vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__clkbuf_2
Xfanout272 net273 vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_31_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13941_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[8\] _03814_ vssd1
+ vssd1 vccd1 vccd1 _03815_ sky130_fd_sc_hd__xor2_1
Xfanout283 net285 vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__buf_2
Xfanout294 net297 vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__buf_2
XANTENNA__08030__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[19\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16660_ clknet_leaf_111_wb_clk_i _02290_ _00356_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_13872_ net1526 net983 _03772_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[7\]
+ sky130_fd_sc_hd__o21a_1
X_15611_ net1149 vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1082 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12823_ net328 net2189 net486 vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__mux2_1
X_16591_ clknet_leaf_134_wb_clk_i _02221_ _00287_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13082__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18330_ net1319 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
XANTENNA__10078__B1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_141_Right_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15542_ net1139 vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12754_ net313 net2337 net495 vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__mux2_1
XANTENNA__09483__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11705_ net548 net356 vssd1 vssd1 vccd1 vccd1 _07517_ sky130_fd_sc_hd__nor2_1
X_18261_ clknet_leaf_37_wb_clk_i _03490_ _01956_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[15\]
+ sky130_fd_sc_hd__dfrtp_4
X_15473_ net1171 vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__inv_2
XANTENNA__11290__A2 _07106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12685_ net2943 net341 vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08691__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_144_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_144_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_84_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17212_ clknet_leaf_154_wb_clk_i _02842_ _00908_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13567__A1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11636_ _04166_ team_05_WB.instance_to_wrap.wishbone.prev_BUSY_O net990 vssd1 vssd1
+ vccd1 vccd1 _07483_ sky130_fd_sc_hd__and3_1
X_14424_ net1207 vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__inv_2
X_18192_ clknet_leaf_41_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[13\]
+ _01887_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09235__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17143_ clknet_leaf_147_wb_clk_i _02773_ _00839_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11567_ net88 net1007 _07354_ _07456_ vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__a22o_1
XANTENNA__12426__S net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11042__A2 _06847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10294__X _06317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08443__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14355_ _04077_ _04127_ _04070_ vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_141_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08994__A1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10518_ _06064_ _06525_ _06529_ vssd1 vssd1 vccd1 vccd1 _06530_ sky130_fd_sc_hd__a21oi_1
X_13306_ net2560 net246 net429 vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__mux2_1
X_14286_ _06369_ _04059_ _06408_ _06387_ vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__or4b_1
XFILLER_0_123_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17074_ clknet_leaf_125_wb_clk_i _02704_ _00770_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold709 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net2123 sky130_fd_sc_hd__dlygate4sd3_1
X_11498_ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[27\] _07408_ net1002
+ vssd1 vssd1 vccd1 vccd1 _07409_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13237_ net234 net2398 net438 vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16025_ net1284 vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__inv_2
X_10449_ _04970_ _05838_ vssd1 vssd1 vccd1 vccd1 _06464_ sky130_fd_sc_hd__xor2_4
XTAP_TAPCELL_ROW_55_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13168_ net236 net2408 net443 vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__mux2_1
XANTENNA__10553__A1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13257__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12119_ _07927_ _07930_ vssd1 vssd1 vccd1 vccd1 _07931_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_72_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09307__Y team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17976_ clknet_leaf_105_wb_clk_i _03315_ _01672_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__dfrtp_1
X_13099_ net224 net2372 net450 vssd1 vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__mux2_1
Xhold1409 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2823 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_144_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14295__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[26\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16927_ clknet_leaf_155_wb_clk_i _02557_ _00623_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_16858_ clknet_leaf_12_wb_clk_i _02488_ _00554_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_140_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15809_ net1277 vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16789_ clknet_leaf_117_wb_clk_i _02419_ _00485_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11505__S net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09330_ _05351_ _05374_ vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_46_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_153_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10188__Y _06215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09474__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09261_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[9\]
+ net834 net830 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__a22o_1
XANTENNA__11281__A2 _07104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08212_ net878 net874 net862 vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__and3_1
XANTENNA__13558__A1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11018__C1 _04170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09192_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[10\]
+ net703 net655 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[10\]
+ _05240_ vssd1 vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08143_ _04220_ _04225_ _04227_ vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__and3b_1
XFILLER_0_43_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout219_A net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08074_ net1027 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[24\]
+ net974 _04186_ vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_116_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload130 clknet_leaf_140_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload130/Y sky130_fd_sc_hd__inv_6
Xclkload141 clknet_leaf_124_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload141/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload152 clknet_leaf_137_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload152/X sky130_fd_sc_hd__clkbuf_4
Xclkload163 clknet_leaf_79_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload163/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_168_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload174 clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload174/Y sky130_fd_sc_hd__inv_8
Xclkload185 clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload185/Y sky130_fd_sc_hd__inv_8
XFILLER_0_141_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1030_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout490_A _03700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13167__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[10\]
+ vssd1 vssd1 vccd1 vccd1 net1428 sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[15\]
+ net818 net790 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__a22o_1
Xhold25 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[22\]
+ vssd1 vssd1 vccd1 vccd1 net1439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[30\] vssd1 vssd1
+ vccd1 vccd1 net1450 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[1\] vssd1 vssd1
+ vccd1 vccd1 net1461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[24\]
+ vssd1 vssd1 vccd1 vccd1 net1472 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_85_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold69 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[11\]
+ vssd1 vssd1 vccd1 vccd1 net1483 sky130_fd_sc_hd__dlygate4sd3_1
X_18387__1369 vssd1 vssd1 vccd1 vccd1 _18387__1369/HI net1369 sky130_fd_sc_hd__conb_1
XFILLER_0_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout922_A _05213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09528_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[3\]
+ net814 _05563_ vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout710_X net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09459_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[5\]
+ net773 net747 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[5\]
+ _05494_ vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__a221o_1
XANTENNA__11272__A2 _07096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08673__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout808_X net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13630__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11009__C1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12470_ net1662 _07836_ _03670_ vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10480__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11421_ _07323_ _07339_ vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08425__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14140_ team_05_WB.instance_to_wrap.CPU_DAT_O\[23\] net504 net912 vssd1 vssd1 vccd1
+ vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[23\] sky130_fd_sc_hd__and3_1
X_11352_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[5\] net508 net359
+ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[1\] vssd1 vssd1 vccd1
+ vccd1 _03388_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08025__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[31\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10303_ net370 _06324_ vssd1 vssd1 vccd1 vccd1 _06325_ sky130_fd_sc_hd__or2_1
X_14071_ _03933_ _03937_ vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__or2_1
X_11283_ _07228_ _07229_ _07243_ vssd1 vssd1 vccd1 vccd1 _07244_ sky130_fd_sc_hd__or3_1
XFILLER_0_120_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13022_ net316 net2822 net463 vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__mux2_1
XANTENNA_input51_A wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10234_ _06068_ _06074_ vssd1 vssd1 vccd1 vccd1 _06259_ sky130_fd_sc_hd__nor2_1
XANTENNA__10535__A1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08312__X _04394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1001 _07345_ vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13077__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1012 _07343_ vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__buf_4
X_17830_ clknet_leaf_76_wb_clk_i _03173_ _01526_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[76\]
+ sky130_fd_sc_hd__dfrtp_1
X_10165_ _06190_ _06191_ _05634_ vssd1 vssd1 vccd1 vccd1 _06192_ sky130_fd_sc_hd__mux2_1
Xfanout1023 net1026 vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__clkbuf_2
Xfanout1034 net1035 vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_50_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1045 net1047 vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__buf_2
Xfanout1056 net1065 vssd1 vssd1 vccd1 vccd1 net1056 sky130_fd_sc_hd__buf_4
X_17761_ clknet_leaf_100_wb_clk_i _03104_ _01457_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14973_ net1087 vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__inv_2
Xfanout1067 net1069 vssd1 vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__buf_4
X_10096_ _06119_ _06122_ net512 vssd1 vssd1 vccd1 vccd1 _06124_ sky130_fd_sc_hd__mux2_1
Xfanout1078 net1108 vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__buf_2
Xfanout1089 net1094 vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__buf_4
XFILLER_0_57_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16712_ clknet_leaf_204_wb_clk_i _02342_ _00408_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13924_ team_05_WB.instance_to_wrap.CPU_DAT_O\[0\] net506 _03799_ vssd1 vssd1 vccd1
+ vccd1 _03800_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17692_ clknet_leaf_86_wb_clk_i _03035_ _01388_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[66\]
+ sky130_fd_sc_hd__dfrtp_1
X_16643_ clknet_leaf_198_wb_clk_i _02273_ _00339_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13855_ team_05_WB.instance_to_wrap.total_design.core.data_mem.last_read net1050
+ vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_18_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12806_ net249 net2385 net486 vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__mux2_1
X_16574_ clknet_leaf_170_wb_clk_i _02204_ _00270_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13786_ _03751_ _03753_ _03756_ _03758_ vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__or4_2
X_10998_ net1045 _06568_ _06975_ net959 vssd1 vssd1 vccd1 vccd1 _06976_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_48_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09456__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18313_ net1405 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
X_15525_ net1170 vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__inv_2
XANTENNA__11263__A2 _07125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12460__A1 _03664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12737_ net226 net2107 net494 vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__mux2_1
XANTENNA__08664__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13540__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18244_ clknet_leaf_59_wb_clk_i net1476 _01939_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15456_ net1155 vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__inv_2
X_12668_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[21\]
+ net341 vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12664__B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14407_ net1523 vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18175_ clknet_leaf_45_wb_clk_i _03474_ _01870_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.key_counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11015__A2 _06609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08416__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11619_ net1612 net1009 net344 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__a22o_1
XANTENNA__12009__X _07821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15387_ net1100 vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__inv_2
XANTENNA__10465__A net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12599_ _03604_ net1813 net203 vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__mux2_1
XANTENNA__09676__D net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17126_ clknet_leaf_117_wb_clk_i _02756_ _00822_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14338_ _05351_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[8\]
+ _04108_ _04109_ _04110_ vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__o2111a_1
Xhold506 net161 vssd1 vssd1 vccd1 vccd1 net1920 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold517 _03300_ vssd1 vssd1 vccd1 vccd1 net1931 sky130_fd_sc_hd__dlygate4sd3_1
Xhold528 team_05_WB.instance_to_wrap.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 net1942
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17057_ clknet_leaf_148_wb_clk_i _02687_ _00753_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold539 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 net1953 sky130_fd_sc_hd__dlygate4sd3_1
X_14269_ team_05_WB.instance_to_wrap.total_design.keypad0.counter\[0\] team_05_WB.instance_to_wrap.total_design.keypad0.counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16152__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16008_ net1112 vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_111_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08222__X _04305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08830_ _04884_ _04885_ _04888_ _04898_ vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__or4_1
Xhold1206 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net2620 sky130_fd_sc_hd__dlygate4sd3_1
X_08761_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[21\]
+ net827 net772 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__a22o_1
Xhold1217 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2631 sky130_fd_sc_hd__dlygate4sd3_1
X_17959_ clknet_leaf_107_wb_clk_i net1880 _01655_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__dfrtp_1
Xhold1228 net136 vssd1 vssd1 vccd1 vccd1 net2642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1239 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net2653 sky130_fd_sc_hd__dlygate4sd3_1
X_08692_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[22\]
+ net641 net612 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[22\]
+ _04764_ vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__a221o_1
XANTENNA__09695__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13228__A0 _06766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_169_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_71_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09447__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09313_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[8\]
+ net753 net750 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__a22o_1
XANTENNA__12451__A1 _03610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11254__A2 _07113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10927__X _06918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13450__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09244_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[9\]
+ net670 net638 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[9\]
+ _05294_ vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1078_A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11006__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09175_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[11\]
+ net798 _05228_ net853 vssd1 vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__a211o_1
XFILLER_0_69_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08407__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09586__D net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1245_A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08126_ _04211_ team_05_WB.instance_to_wrap.total_design.keypad0.next_rows\[1\] vssd1
+ vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09080__B1 _04417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08057_ team_05_WB.instance_to_wrap.total_design.core.data_mem.state\[1\] vssd1 vssd1
+ vccd1 vccd1 _04177_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1033_X net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout493_X net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout872_A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08959_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[15\]
+ net687 net640 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout660_X net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout758_X net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11493__X _07404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11970_ _07528_ _07781_ vssd1 vssd1 vccd1 vccd1 _07782_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_16_Left_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10921_ _06784_ _06785_ _06787_ _06879_ vssd1 vssd1 vccd1 vccd1 _06913_ sky130_fd_sc_hd__a211o_1
XFILLER_0_86_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout925_X net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10852_ _06847_ _06848_ _06834_ vssd1 vssd1 vccd1 vccd1 _06849_ sky130_fd_sc_hd__a21bo_1
X_13640_ net2791 net260 net389 vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09438__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11245__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10783_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[28\] net1040 vssd1
+ vssd1 vccd1 vccd1 _06780_ sky130_fd_sc_hd__or2_1
XANTENNA__12442__A1 _03661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13571_ net2027 net253 net396 vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__mux2_1
XANTENNA__08646__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14309__X _04082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13360__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08110__A2 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15310_ net1188 vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__inv_2
X_12522_ net1621 _03620_ net208 vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__mux2_1
X_16290_ net1165 vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_23_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15241_ net1221 vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__inv_2
X_12453_ net1615 _03620_ net212 vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11404_ net2154 _07329_ vssd1 vssd1 vccd1 vccd1 _07333_ sky130_fd_sc_hd__nor2_1
X_12384_ net1627 _03645_ _03660_ vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__mux2_1
X_15172_ net1229 vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__inv_2
XANTENNA__09071__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11335_ _07292_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.next_rows\[3\]
+ sky130_fd_sc_hd__inv_2
X_14123_ _03985_ _03986_ vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12704__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14054_ _03921_ _03922_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__and2_1
X_11266_ net2440 net732 _07211_ _07227_ vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__o22a_1
XANTENNA__09374__A1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10217_ _06221_ _06241_ _06242_ net537 vssd1 vssd1 vccd1 vccd1 _06243_ sky130_fd_sc_hd__a31o_1
X_13005_ net226 net2588 net463 vssd1 vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__mux2_1
X_11197_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[70\] _07128_
+ _07129_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[62\] vssd1 vssd1
+ vccd1 vccd1 _07162_ sky130_fd_sc_hd__a22o_1
XANTENNA__08202__B net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17813_ clknet_leaf_103_wb_clk_i _03156_ _01509_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[123\]
+ sky130_fd_sc_hd__dfrtp_1
X_10148_ net520 _06175_ _06172_ net531 vssd1 vssd1 vccd1 vccd1 _06176_ sky130_fd_sc_hd__o211a_1
XANTENNA__13535__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11844__A _07623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17744_ clknet_leaf_94_wb_clk_i _03087_ _01440_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10079_ net2268 net197 net540 vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__mux2_1
X_14956_ net1071 vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_89_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12659__B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13907_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[25\]
+ net559 net575 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[25\]
+ net986 vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__a221o_1
X_17675_ clknet_leaf_75_wb_clk_i _03018_ _01371_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[113\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08885__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14887_ net1176 vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10692__B1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16626_ clknet_leaf_133_wb_clk_i _02256_ _00322_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13838_ net1519 net578 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[16\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_134_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09429__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11236__A2 _07120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12433__A1 _07816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16557_ clknet_leaf_161_wb_clk_i _02187_ _00253_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08637__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13769_ _03738_ _03739_ _03741_ vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__or3_1
XANTENNA__13270__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15508_ net1172 vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_21_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16488_ clknet_leaf_201_wb_clk_i _02118_ _00184_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_135_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18227_ clknet_leaf_62_wb_clk_i net1498 _01922_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15439_ net1253 vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12962__X _03710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09984__A net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18158_ clknet_leaf_138_wb_clk_i _03461_ _01854_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_152_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09062__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold303 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[36\] vssd1 vssd1
+ vccd1 vccd1 net1717 sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[71\] vssd1 vssd1
+ vccd1 vccd1 net1728 sky130_fd_sc_hd__dlygate4sd3_1
X_17109_ clknet_leaf_175_wb_clk_i _02739_ _00805_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold325 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[32\] vssd1 vssd1
+ vccd1 vccd1 net1739 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12614__S net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18089_ clknet_leaf_79_wb_clk_i _03412_ _01785_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[6\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold336 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[3\]
+ vssd1 vssd1 vccd1 vccd1 net1750 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold347 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[26\] vssd1 vssd1
+ vccd1 vccd1 net1761 sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[58\] vssd1 vssd1
+ vccd1 vccd1 net1772 sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[98\] vssd1 vssd1
+ vccd1 vccd1 net1783 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ _05285_ _05817_ _05957_ _05938_ _05824_ vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__a311o_1
XFILLER_0_111_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout805 _04393_ vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__buf_4
Xfanout816 _04388_ vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_68_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09862_ _04799_ _05888_ _05889_ vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__and3_1
Xfanout827 net828 vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__buf_4
Xfanout838 net840 vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout849 _04370_ vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__clkbuf_8
Xhold1003 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2417 sky130_fd_sc_hd__dlygate4sd3_1
X_08813_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[18\]
+ net617 net610 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__a22o_1
X_09793_ _05823_ vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__inv_2
Xhold1014 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2428 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1025 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1036 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2450 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13445__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1047 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 net2461 sky130_fd_sc_hd__dlygate4sd3_1
X_08744_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[21\]
+ net684 net649 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[21\]
+ _04800_ vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__a221o_1
Xhold1058 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net2472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1069 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 net2483 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08325__C1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08675_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[23\]
+ net838 net779 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[23\]
+ _04748_ vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout453_A _03713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12424__A1 _03663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11227__A2 _07096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08628__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13180__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout339_X net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout718_A _04286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10435__A0 _06284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09840__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18045__Q team_05_WB.instance_to_wrap.total_design.data_from_keypad\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09227_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[10\]
+ net590 _05269_ _05278_ vssd1 vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_63_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09158_ net1022 _04231_ _04241_ vssd1 vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__or3_4
XANTENNA__09894__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[14\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09053__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08109_ net1029 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__and2b_1
XFILLER_0_121_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12524__S net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09089_ _05145_ vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__inv_2
XANTENNA__08800__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11120_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[5\] _07037_
+ _07070_ vssd1 vssd1 vccd1 vccd1 _07087_ sky130_fd_sc_hd__o21a_4
XANTENNA__13688__A0 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold870 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 net2284 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout875_X net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold881 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2295 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11051_ _06837_ _06843_ _06842_ vssd1 vssd1 vccd1 vccd1 _07019_ sky130_fd_sc_hd__a21o_1
Xhold892 team_05_WB.instance_to_wrap.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 net2306
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10002_ _06027_ _06030_ net513 vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__mux2_1
XANTENNA__13355__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14810_ net1056 vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__inv_2
X_15790_ net1297 vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09659__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14741_ net1079 vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__inv_2
XANTENNA_input14_A DAT_I[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11953_ _07737_ _07750_ _07762_ _07764_ vssd1 vssd1 vccd1 vccd1 _07765_ sky130_fd_sc_hd__a22oi_4
XANTENNA__08867__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08331__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17460_ clknet_leaf_56_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[28\]
+ _01156_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10904_ net1044 net957 vssd1 vssd1 vccd1 vccd1 _06899_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_28_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14672_ net1182 vssd1 vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__inv_2
X_11884_ _07652_ _07660_ vssd1 vssd1 vccd1 vccd1 _07696_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_84_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16411_ clknet_leaf_189_wb_clk_i _02041_ _00107_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13623_ net1952 net327 net393 vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17391_ clknet_leaf_58_wb_clk_i net1442 _01087_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10835_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[5\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06832_ sky130_fd_sc_hd__nand2_1
XANTENNA__08619__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13090__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16342_ net1131 vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__inv_2
X_13554_ net2093 net330 net402 vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09292__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10766_ _06492_ net347 _06758_ _06763_ vssd1 vssd1 vccd1 vccd1 _06764_ sky130_fd_sc_hd__o211a_1
XANTENNA__09831__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12505_ net1783 _07836_ _03673_ vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16273_ net1119 vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__inv_2
X_10697_ net369 net348 _06698_ _06695_ vssd1 vssd1 vccd1 vccd1 _06699_ sky130_fd_sc_hd__o31a_1
X_13485_ net304 net2264 net410 vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__mux2_1
X_18012_ clknet_leaf_82_wb_clk_i _03351_ _01708_ vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__dfrtp_1
X_15224_ net1244 vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__inv_2
X_12436_ _03641_ net1901 net214 vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08398__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15155_ net1212 vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__inv_2
XANTENNA__12434__S _03668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12367_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[30\] net996 _03626_
+ net545 vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__a211o_2
XFILLER_0_2_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14106_ _03952_ _03964_ vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__nand2_1
XANTENNA__11558__B _07452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11318_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[40\] _07091_
+ _07127_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[120\] _07266_
+ vssd1 vssd1 vccd1 vccd1 _07277_ sky130_fd_sc_hd__a221o_1
X_12298_ _03569_ _03575_ _03557_ vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__a21bo_1
X_15086_ net1180 vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_39_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14340__A1 _05208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14037_ _03877_ _03879_ _03906_ vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__a21o_1
X_11249_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[3\] _07100_ _07169_
+ _07208_ _07210_ vssd1 vssd1 vccd1 vccd1 _07211_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_129_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14340__B2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12351__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11845__Y _07657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13265__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15988_ net1129 vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1068 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17727_ clknet_leaf_86_wb_clk_i _03070_ _01423_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09044__A _05078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14939_ net1098 vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08460_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[28\]
+ net784 net773 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[28\]
+ _04538_ vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__a221o_1
X_17658_ clknet_leaf_92_wb_clk_i _03001_ _01354_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[96\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16609_ clknet_leaf_150_wb_clk_i _02239_ _00305_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11209__A2 _07109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08391_ _04470_ vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__inv_2
XFILLER_0_147_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12609__S net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17589_ clknet_leaf_73_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[26\]
+ _01285_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_102_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10918__A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11513__S net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09283__B1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09822__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09012_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[14\]
+ net689 net599 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_171_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_171_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09035__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold100 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[25\] vssd1 vssd1
+ vccd1 vccd1 net1514 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold111 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[18\]
+ vssd1 vssd1 vccd1 vccd1 net1525 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout201_A _03683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold122 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[31\]
+ vssd1 vssd1 vccd1 vccd1 net1536 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12590__A0 _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold133 team_05_WB.instance_to_wrap.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 net1547
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[20\]
+ vssd1 vssd1 vccd1 vccd1 net1558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[22\]
+ vssd1 vssd1 vccd1 vccd1 net1569 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[3\]
+ vssd1 vssd1 vccd1 vccd1 net1580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 net80 vssd1 vssd1 vccd1 vccd1 net1591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[7\]
+ vssd1 vssd1 vccd1 vccd1 net1602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[24\]
+ vssd1 vssd1 vccd1 vccd1 net1613 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout602 net605 vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__clkbuf_8
X_09914_ net525 net523 vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__nor2_1
Xfanout613 _04319_ vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__buf_4
XFILLER_0_0_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout624 _04316_ vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1110_A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout635 _04313_ vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__buf_4
Xfanout646 net647 vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__buf_4
XANTENNA_input6_A DAT_I[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09845_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[20\]
+ net794 net790 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__a22o_1
Xfanout657 net659 vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout570_A _04344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11696__A2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[17\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout668 net671 vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08410__X _04490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout679 _04302_ vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout289_X net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout668_A net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13175__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13028__X _03712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09776_ _05804_ _05806_ _05597_ vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_126_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ _04777_ _04797_ vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout456_X net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout835_A net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[23\]
+ net634 net595 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[23\]
+ _04718_ vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_1_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout623_X net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12519__S net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08589_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[25\]
+ net773 net743 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[25\]
+ _04664_ vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10620_ _06048_ _06328_ vssd1 vssd1 vccd1 vccd1 _06626_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09813__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10551_ _06490_ _06560_ net528 vssd1 vssd1 vccd1 vccd1 _06561_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11620__A2 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10482_ _06094_ _06495_ vssd1 vssd1 vccd1 vccd1 _06496_ sky130_fd_sc_hd__or2_1
X_13270_ net234 net2426 net435 vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__mux2_1
XANTENNA__09026__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12221_ _08010_ _08021_ _03512_ _03515_ vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_103_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12581__A0 _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08785__C1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12152_ _07950_ _07954_ _07960_ _07952_ vssd1 vssd1 vccd1 vccd1 _07964_ sky130_fd_sc_hd__o22ai_2
X_11103_ _04161_ _04162_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[3\]
+ _07061_ vssd1 vssd1 vccd1 vccd1 _07070_ sky130_fd_sc_hd__or4b_2
XFILLER_0_20_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_169_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_169_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10850__X _06847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16960_ clknet_leaf_132_wb_clk_i _02590_ _00656_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_12083_ _07894_ vssd1 vssd1 vccd1 vccd1 _07895_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15911_ net1291 vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__inv_2
X_11034_ _06832_ _06833_ _06849_ vssd1 vssd1 vccd1 vccd1 _07005_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16891_ clknet_leaf_191_wb_clk_i _02521_ _00587_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13085__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08552__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15842_ net1296 vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_34_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11439__A2 _07351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15773_ net1290 vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__inv_2
X_12985_ net300 net2340 net466 vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__mux2_1
X_17512_ clknet_leaf_113_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[15\]
+ _01208_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08304__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14724_ net1229 vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__inv_2
X_11936_ _07722_ _07724_ _07745_ _07747_ vssd1 vssd1 vccd1 vccd1 _07748_ sky130_fd_sc_hd__or4_1
XFILLER_0_86_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17443_ clknet_leaf_65_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[11\]
+ _01139_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_14655_ net1178 vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__inv_2
XANTENNA__12429__S net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11867_ _07648_ _07678_ vssd1 vssd1 vccd1 vccd1 _07679_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13606_ net2591 net263 net392 vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17374_ clknet_leaf_79_wb_clk_i net1421 _01070_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10818_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[13\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06815_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_60_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14586_ net1056 vssd1 vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11798_ _07607_ _07609_ vssd1 vssd1 vccd1 vccd1 _07610_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16325_ net1116 vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13537_ net2020 net247 net400 vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10749_ net525 _06679_ net335 vssd1 vssd1 vccd1 vccd1 _06748_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_131_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16256_ net1138 vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__inv_2
X_13468_ net235 net2455 net410 vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__mux2_1
XANTENNA__12672__B net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15207_ net1202 vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__inv_2
X_12419_ _03614_ net1868 net214 vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__mux2_1
X_16187_ net1135 vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__inv_2
XANTENNA__11375__A1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13399_ net2069 net225 net418 vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__mux2_1
XANTENNA__09684__D net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15138_ net1228 vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_58_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08791__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15069_ net1092 vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__inv_2
XANTENNA__09326__X team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08230__X _04313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_155_Right_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08543__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09630_ _05654_ _05655_ _05656_ _05657_ vssd1 vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__or4_1
XFILLER_0_156_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09561_ _04149_ net955 _04268_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_104_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11591__X _07472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10638__B1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08512_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[27\]
+ net851 net842 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[27\]
+ _04589_ vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__a221o_1
X_09492_ net573 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[4\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[4\] vssd1 vssd1 vccd1
+ vccd1 _05531_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_19_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_121_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08443_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[28\]
+ net650 net603 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[28\]
+ _04517_ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_173_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08374_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[30\]
+ net819 net807 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[30\]
+ _04454_ vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__a221o_1
XFILLER_0_147_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout416_A _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1158_A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09008__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout204_X net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11366__A1 team_05_WB.instance_to_wrap.total_design.data_from_keypad\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08782__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14304__A1 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14304__B2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[30\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12802__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout410 _03728_ vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout421 net422 vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__clkbuf_8
Xfanout432 _03722_ vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__buf_6
Xfanout443 _03716_ vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__buf_4
Xfanout454 _03713_ vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__buf_6
XANTENNA_fanout573_X net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout465 _03710_ vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14302__B _04552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08534__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout476 net479 vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__buf_6
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09828_ _05845_ _05847_ _05849_ _05858_ vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__or4_1
Xfanout487 _03703_ vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__buf_4
Xfanout498 net499 vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__buf_4
XANTENNA__08300__B net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12618__A1 _07791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout740_X net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09759_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[0\]
+ net647 net610 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout838_X net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13633__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12770_ net226 net2710 net489 vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09495__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11721_ _07519_ _07525_ vssd1 vssd1 vccd1 vccd1 _07533_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_81_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10644__A3 _06049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14440_ net1218 vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__inv_2
XFILLER_0_167_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11652_ net10 net991 net918 team_05_WB.instance_to_wrap.CPU_DAT_O\[17\] vssd1 vssd1
+ vccd1 vccd1 _03276_ sky130_fd_sc_hd__a22o_1
XANTENNA__09247__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08028__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[21\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10603_ net890 _06609_ _06608_ net555 vssd1 vssd1 vccd1 vccd1 _06610_ sky130_fd_sc_hd__a211o_1
XFILLER_0_119_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14371_ _04143_ _06002_ _04123_ vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__mux2_1
X_11583_ net1988 net1005 _07376_ net357 vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16110_ net1152 vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__inv_2
X_13322_ net2018 net314 net430 vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17090_ clknet_leaf_16_wb_clk_i _02720_ _00786_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10534_ _06468_ _06544_ net529 vssd1 vssd1 vccd1 vccd1 _06545_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16041_ net1287 vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__inv_2
X_13253_ net294 net2166 net439 vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__mux2_1
X_10465_ net382 _06479_ vssd1 vssd1 vccd1 vccd1 _06480_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12554__A0 _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12204_ _08015_ vssd1 vssd1 vccd1 vccd1 _08016_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10396_ _05881_ _06051_ _06055_ _05884_ vssd1 vssd1 vccd1 vccd1 _06414_ sky130_fd_sc_hd__o2bb2a_1
X_13184_ net295 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[8\]
+ net443 vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12135_ _07943_ _07946_ vssd1 vssd1 vccd1 vccd1 _07947_ sky130_fd_sc_hd__nand2_1
XANTENNA__08773__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17992_ clknet_leaf_83_wb_clk_i _03331_ _01688_ vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12712__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16943_ clknet_leaf_135_wb_clk_i _02573_ _00639_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_12066_ _07865_ _07877_ vssd1 vssd1 vccd1 vccd1 _07878_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_53_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Left_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08525__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11017_ _06827_ _06853_ _06852_ vssd1 vssd1 vccd1 vccd1 _06991_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10232__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16874_ clknet_leaf_181_wb_clk_i _02504_ _00570_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1032 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08210__B net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15825_ net1267 vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13543__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15324__A net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15756_ net1300 vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12968_ net242 net2162 net467 vssd1 vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_66_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_36_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12667__B net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14707_ net1213 vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__inv_2
XANTENNA__11293__B1 _07103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11919_ _07692_ _07698_ _07694_ _07688_ vssd1 vssd1 vccd1 vccd1 _07731_ sky130_fd_sc_hd__a2bb2o_1
X_15687_ net1160 vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12899_ net222 net2808 net474 vssd1 vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17426_ clknet_leaf_56_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[26\]
+ _01122_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14638_ net1187 vssd1 vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09238__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17357_ clknet_leaf_35_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[21\]
+ _01053_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14569_ net1222 vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11596__A1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16308_ net1160 vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__inv_2
XFILLER_0_166_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08090_ net1023 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[16\]
+ net970 _04194_ vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17288_ clknet_leaf_204_wb_clk_i _02918_ _00984_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload20 clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload20/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_67_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16239_ net1135 vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload31 clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload31/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload42 clknet_leaf_191_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload42/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__12545__A0 _07857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload53 clknet_leaf_176_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload53/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_24_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload64 clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload64/Y sky130_fd_sc_hd__inv_12
XTAP_TAPCELL_ROW_77_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload75 clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload75/Y sky130_fd_sc_hd__inv_8
XFILLER_0_140_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire374_X net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09992__A net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload86 clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload86/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09410__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload97 clknet_leaf_59_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload97/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__17982__Q net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12622__S net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08992_ _05047_ _05049_ _05051_ _05053_ vssd1 vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_166_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_75_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11520__A1 _07346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10323__A2 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08921__C1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09613_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[2\]
+ net877 net865 net861 vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_123_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13453__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout366_A net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09544_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[3\]
+ net699 net606 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__a22o_1
XANTENNA__09477__B1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09475_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[4\]
+ net838 net779 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08426_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[29\]
+ net831 net791 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[29\]
+ _04499_ vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__a221o_1
XFILLER_0_136_616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09229__B1 _05260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08357_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[30\]
+ net670 net616 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[30\]
+ _04437_ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout700_A _04293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11587__A1 _07354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload3 clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload3/Y sky130_fd_sc_hd__inv_6
XFILLER_0_19_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1063_X net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout419_X net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08288_ net949 net938 net935 vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__and3_4
XFILLER_0_150_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18280__A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12536__A0 _07821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10250_ net893 _06273_ vssd1 vssd1 vccd1 vccd1 _06274_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09401__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout690_X net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11496__X _07407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout788_X net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08755__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13628__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10181_ _06012_ _06023_ net516 vssd1 vssd1 vccd1 vccd1 _06208_ sky130_fd_sc_hd__mux2_1
XANTENNA__12532__S _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14313__A _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1205 net1206 vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__buf_2
Xfanout1216 net1217 vssd1 vssd1 vccd1 vccd1 net1216 sky130_fd_sc_hd__buf_4
Xfanout1227 net1234 vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__buf_2
XANTENNA__08311__A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout240 net241 vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__buf_2
Xfanout1238 net1240 vssd1 vssd1 vccd1 vccd1 net1238 sky130_fd_sc_hd__buf_4
Xfanout1249 net1252 vssd1 vssd1 vccd1 vccd1 net1249 sky130_fd_sc_hd__buf_4
XANTENNA__09704__A1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[20\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08507__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout262 _06480_ vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__clkbuf_2
X_13940_ _03812_ _03813_ vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__nand2_1
XANTENNA__09704__B2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout273 _06518_ vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_31_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout284 net285 vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout295 net297 vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09180__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13871_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[7\]
+ net559 net575 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[7\]
+ net986 vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__a221o_1
X_15610_ net1168 vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__inv_2
XANTENNA__11672__A team_05_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13363__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12822_ net313 net2586 net487 vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__mux2_1
X_16590_ clknet_leaf_172_wb_clk_i _02220_ _00286_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11275__B1 _07116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15541_ net1133 vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12753_ net318 net2387 net493 vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11704_ net501 vssd1 vssd1 vccd1 vccd1 _07516_ sky130_fd_sc_hd__inv_2
X_18260_ clknet_leaf_33_wb_clk_i _03489_ _01955_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[14\]
+ sky130_fd_sc_hd__dfrtp_4
X_15472_ net1166 vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__inv_2
X_12684_ net2813 net342 vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__and2_1
XFILLER_0_139_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17211_ clknet_leaf_191_wb_clk_i _02841_ _00907_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_14423_ net1104 vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__inv_2
X_11635_ team_05_WB.instance_to_wrap.wishbone.curr_state\[1\] net1 vssd1 vssd1 vccd1
+ vccd1 _07482_ sky130_fd_sc_hd__nand2_1
X_18191_ clknet_leaf_40_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[12\]
+ _01886_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12707__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17142_ clknet_leaf_151_wb_clk_i _02772_ _00838_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14354_ _04125_ _04126_ _04073_ _04074_ vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__a211o_1
X_11566_ net1780 net1007 net727 _07402_ vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_184_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_184_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13305_ net2084 net228 net430 vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__mux2_1
X_10517_ _05104_ _06056_ _06160_ _06509_ _06528_ vssd1 vssd1 vccd1 vccd1 _06529_ sky130_fd_sc_hd__a221o_1
XANTENNA__08994__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[15\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17073_ clknet_leaf_172_wb_clk_i _02703_ _00769_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_14285_ _06424_ _06445_ _06464_ _04058_ vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__or4b_1
X_11497_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[27\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[27\]
+ net1034 vssd1 vssd1 vccd1 vccd1 _07408_ sky130_fd_sc_hd__mux2_1
XANTENNA__12527__A0 _07812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08205__B net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_113_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_113_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16024_ net1284 vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__inv_2
X_13236_ net239 net2549 net438 vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10448_ _04970_ _05970_ vssd1 vssd1 vccd1 vccd1 _06463_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13538__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08746__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11847__A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12442__S net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13167_ net240 net2871 net442 vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__mux2_1
X_10379_ _06199_ _06397_ net372 vssd1 vssd1 vccd1 vccd1 _06398_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12118_ _07926_ _07929_ _07921_ _07922_ vssd1 vssd1 vccd1 vccd1 _07930_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_72_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17975_ clknet_leaf_106_wb_clk_i _03314_ _01671_ vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__dfrtp_1
X_13098_ net218 net2420 net451 vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_144_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12049_ _07369_ _07468_ _07841_ vssd1 vssd1 vccd1 vccd1 _07861_ sky130_fd_sc_hd__or3_1
X_16926_ clknet_leaf_185_wb_clk_i _02556_ _00622_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09171__A2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16857_ clknet_leaf_10_wb_clk_i _02487_ _00553_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13273__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_159_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_88_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15054__A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15808_ net1276 vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09459__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16788_ clknet_leaf_114_wb_clk_i _02418_ _00484_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15739_ net1301 vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09260_ _05309_ _05310_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[9\]
+ sky130_fd_sc_hd__nand2_1
XANTENNA__08682__A1 _04344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17977__Q net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10613__A2_N net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08211_ _04232_ net962 _04271_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[17\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[18\] vssd1 vssd1
+ vccd1 vccd1 _04294_ sky130_fd_sc_hd__o311a_1
X_17409_ clknet_leaf_65_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[9\]
+ _01105_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_09191_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[10\]
+ net700 net636 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[10\]
+ _05243_ vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__a221o_1
X_18389_ net913 vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12617__S _03682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10485__X _06499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12766__A0 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11569__B2 _07414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08142_ team_05_WB.instance_to_wrap.total_design.keypad0.key_counter\[0\] _04219_
+ team_05_WB.instance_to_wrap.total_design.keypad0.key_counter\[1\] vssd1 vssd1 vccd1
+ vccd1 _04227_ sky130_fd_sc_hd__a21o_1
X_08073_ net1027 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__and2b_1
XFILLER_0_114_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08985__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload120 clknet_leaf_122_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload120/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_116_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload131 clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload131/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_116_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload142 clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload142/Y sky130_fd_sc_hd__bufinv_16
Xclkload153 clknet_leaf_71_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload153/Y sky130_fd_sc_hd__inv_12
Xclkload164 clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload164/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_114_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload175 clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload175/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_168_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload186 clknet_leaf_95_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload186/Y sky130_fd_sc_hd__inv_6
Xmax_cap952 _04278_ vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__buf_1
XANTENNA__08198__B1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[19\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13448__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08737__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_198_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08975_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[15\]
+ net829 net810 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__a22o_1
Xhold15 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[19\]
+ vssd1 vssd1 vccd1 vccd1 net1429 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout483_A _03704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold26 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[0\]
+ vssd1 vssd1 vccd1 vccd1 net1440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[5\]
+ vssd1 vssd1 vccd1 vccd1 net1451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[20\] vssd1 vssd1
+ vccd1 vccd1 net1462 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09698__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold59 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09162__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1071 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout650_A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08370__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13183__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout748_A net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11257__B1 _07108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09527_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[3\]
+ net850 net794 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[3\]
+ _05564_ vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout915_A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout536_X net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1278_X net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09458_ _05496_ _05497_ _05498_ _05499_ vssd1 vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__or4_1
XFILLER_0_94_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08409_ _04474_ _04486_ _04487_ _04488_ vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__or4_1
XFILLER_0_109_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12527__S _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09389_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[6\]
+ net680 net649 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout703_X net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11420_ net2117 _07322_ vssd1 vssd1 vccd1 vccd1 _07339_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11351_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[6\] net508 net359
+ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[2\] vssd1 vssd1 vccd1
+ vccd1 _03389_ sky130_fd_sc_hd__a22o_1
XANTENNA__08976__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10302_ net526 _06222_ vssd1 vssd1 vccd1 vccd1 _06324_ sky130_fd_sc_hd__nand2_1
X_14070_ _03933_ _03937_ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_89_Left_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11282_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[82\] _07126_
+ _07127_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[122\] _07242_
+ vssd1 vssd1 vccd1 vccd1 _07243_ sky130_fd_sc_hd__a221o_1
XFILLER_0_131_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13021_ net319 net2564 net462 vssd1 vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__mux2_1
XANTENNA__08728__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13358__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10233_ net1021 _04594_ net553 vssd1 vssd1 vccd1 vccd1 _06258_ sky130_fd_sc_hd__a21oi_1
XANTENNA_input44_A wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1002 _07345_ vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__clkbuf_4
X_10164_ _06042_ _06079_ net521 vssd1 vssd1 vccd1 vccd1 _06191_ sky130_fd_sc_hd__mux2_1
Xfanout1013 net1014 vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__buf_2
Xfanout1024 net1026 vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_50_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1035 net1036 vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1046 net1047 vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__buf_1
X_17760_ clknet_leaf_90_wb_clk_i _03103_ _01456_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1057 net1058 vssd1 vssd1 vccd1 vccd1 net1057 sky130_fd_sc_hd__buf_4
X_14972_ net1083 vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__inv_2
X_10095_ _06122_ vssd1 vssd1 vccd1 vccd1 _06123_ sky130_fd_sc_hd__inv_2
Xfanout1068 net1069 vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__buf_4
Xfanout1079 net1086 vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__buf_4
X_13923_ team_05_WB.instance_to_wrap.total_design.data_from_keypad\[0\] _07451_ vssd1
+ vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__and2_1
XANTENNA__09153__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16711_ clknet_leaf_202_wb_clk_i _02341_ _00407_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17691_ clknet_leaf_90_wb_clk_i _03034_ _01387_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[65\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13093__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16642_ clknet_leaf_8_wb_clk_i _02272_ _00338_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13854_ team_05_WB.instance_to_wrap.total_design.core.data_mem.last_read net1050
+ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_98_Left_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11248__B1 _07127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12805_ net228 net2304 net486 vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__mux2_1
X_16573_ clknet_leaf_131_wb_clk_i _02203_ _00269_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13785_ _03754_ _03755_ _03757_ vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__or3_1
X_10997_ _04170_ _06860_ _06974_ vssd1 vssd1 vccd1 vccd1 _06975_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_48_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15524_ net1170 vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__inv_2
X_18312_ net1404 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
XFILLER_0_69_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12736_ net232 net2698 net494 vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18243_ clknet_leaf_59_wb_clk_i net1450 _01938_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15455_ net1156 vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__inv_2
XANTENNA__12437__S net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12667_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[22\]
+ net342 vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__and2_1
X_14406_ net1539 vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18174_ clknet_leaf_45_wb_clk_i _03473_ _01869_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.key_counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_137_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11618_ net1914 net1009 _07472_ _07478_ vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__a22o_1
X_15386_ net1062 vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__inv_2
X_12598_ _03664_ net1888 net204 vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10759__C1 _06756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17125_ clknet_leaf_178_wb_clk_i _02755_ _00821_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_163_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08967__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14337_ _05035_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[15\]
+ _05078_ _05099_ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__o2bb2a_1
X_11549_ _07414_ _07438_ vssd1 vssd1 vccd1 vccd1 _07460_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold507 team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.next_next_fetch vssd1
+ vssd1 vccd1 vccd1 net1921 sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[23\] vssd1 vssd1
+ vccd1 vccd1 net1932 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold529 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[8\] vssd1 vssd1
+ vccd1 vccd1 net1943 sky130_fd_sc_hd__dlygate4sd3_1
X_17056_ clknet_leaf_129_wb_clk_i _02686_ _00752_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_74_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14268_ _04017_ _04043_ _04047_ vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__nor3_1
XFILLER_0_150_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12680__B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16007_ net1114 vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13268__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08719__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13219_ net303 net2366 net352 vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__mux2_1
XANTENNA__15049__A net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14199_ _04003_ net728 _04002_ vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__and3b_1
XFILLER_0_148_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_111_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09392__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1207 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2621 sky130_fd_sc_hd__dlygate4sd3_1
X_08760_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[21\]
+ net796 net769 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[21\]
+ _04831_ vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__a221o_1
XANTENNA__12900__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1218 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 net2632 sky130_fd_sc_hd__dlygate4sd3_1
X_17958_ clknet_leaf_107_wb_clk_i _03297_ _01654_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_81_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold1229 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2643 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09144__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16909_ clknet_leaf_159_wb_clk_i _02539_ _00605_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_08691_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[22\]
+ net692 net673 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__a22o_1
X_17889_ clknet_leaf_100_wb_clk_i _03232_ _01585_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_10_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08352__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11239__B1 _07129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12987__A0 _06655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09312_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[8\]
+ net808 net743 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[8\]
+ _05359_ vssd1 vssd1 vccd1 vccd1 _05360_ sky130_fd_sc_hd__a221o_1
XANTENNA__15512__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10552__A2_N _06051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10998__C1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09243_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[9\]
+ net685 net595 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18245__D net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout231_A _06367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17500__Q team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout329_A _06705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09174_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[11\]
+ net748 net745 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13400__A1 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08125_ net151 _04212_ net152 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.next_rows\[1\]
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08958__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08056_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[30\] vssd1 vssd1
+ vccd1 vccd1 _04176_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09368__C1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13178__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10517__A2 _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09383__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11190__A2 _07091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout865_A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout486_X net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08591__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08958_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[15\]
+ net707 net636 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[15\]
+ _05020_ vssd1 vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__a221o_1
XANTENNA__12810__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09135__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout653_X net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08889_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[17\]
+ net805 net764 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[17\]
+ _04954_ vssd1 vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__a221o_1
X_10920_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[27\] net566 _06911_
+ _06912_ vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__a22o_1
X_10851_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[4\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06848_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout820_X net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13641__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1090 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13570_ net2056 net247 net398 vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__mux2_1
X_10782_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[28\] net1040 vssd1
+ vssd1 vccd1 vccd1 _06779_ sky130_fd_sc_hd__nand2_1
XANTENNA__09843__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12521_ net1646 _03644_ net209 vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15240_ net1220 vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__inv_2
X_12452_ net1700 _03644_ net213 vssd1 vssd1 vccd1 vccd1 _03181_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08036__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11403_ _07331_ _07332_ vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__and2_1
X_15171_ net1208 vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__inv_2
X_12383_ net1762 _03632_ net217 vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14122_ _03971_ _03974_ _03978_ vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_10_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11334_ net153 net154 net151 net152 vssd1 vssd1 vccd1 vccd1 _07292_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_10_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09419__X team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08157__A_N team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13088__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14053_ _03890_ _03898_ _03920_ vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__or3_1
X_11265_ _07213_ _07216_ _07217_ _07226_ vssd1 vssd1 vccd1 vccd1 _07227_ sky130_fd_sc_hd__or4_1
X_13004_ net232 net2802 net462 vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__mux2_1
XANTENNA__09374__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10216_ net333 _06232_ _06237_ net336 _06233_ vssd1 vssd1 vccd1 vccd1 _06242_ sky130_fd_sc_hd__o221a_1
X_11196_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[22\] _07125_
+ _07130_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[102\] _07149_
+ vssd1 vssd1 vccd1 vccd1 _07161_ sky130_fd_sc_hd__a221o_1
XANTENNA__11181__A2 _07104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08582__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08202__C net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17812_ clknet_leaf_77_wb_clk_i _03155_ _01508_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12720__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10147_ _06173_ _06174_ vssd1 vssd1 vccd1 vccd1 _06175_ sky130_fd_sc_hd__nand2_1
XANTENNA__09126__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17743_ clknet_leaf_86_wb_clk_i _03086_ _01439_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[53\]
+ sky130_fd_sc_hd__dfrtp_1
X_14955_ net1072 vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__inv_2
X_10078_ _06084_ _06106_ net383 vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__o21a_4
XANTENNA__08334__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13906_ net1613 net982 _03789_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[24\]
+ sky130_fd_sc_hd__o21a_1
X_17674_ clknet_leaf_98_wb_clk_i _03017_ _01370_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[112\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08993__X team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[15\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14886_ net1247 vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__inv_2
XFILLER_0_159_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10692__A1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13837_ net1477 net578 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[15\]
+ sky130_fd_sc_hd__and2_1
X_16625_ clknet_leaf_122_wb_clk_i _02255_ _00321_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13551__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16556_ clknet_leaf_0_wb_clk_i _02186_ _00252_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13768_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[29\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[28\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[31\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__or4_1
XFILLER_0_70_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09834__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12675__B net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15507_ net1172 vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_63_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12719_ net313 net2280 net498 vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__mux2_1
X_16487_ clknet_leaf_201_wb_clk_i _02117_ _00183_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13699_ _07480_ _07491_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10995__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15438_ net1258 vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__inv_2
X_18226_ clknet_leaf_68_wb_clk_i net1452 _01921_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_135_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15369_ net1214 vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__inv_2
X_18157_ clknet_leaf_171_wb_clk_i _03460_ _01853_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16163__A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12691__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold304 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[120\] vssd1 vssd1
+ vccd1 vccd1 net1718 sky130_fd_sc_hd__dlygate4sd3_1
X_17108_ clknet_leaf_114_wb_clk_i _02738_ _00804_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold315 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[42\] vssd1 vssd1
+ vccd1 vccd1 net1729 sky130_fd_sc_hd__dlygate4sd3_1
X_18088_ clknet_leaf_79_wb_clk_i _03411_ _01784_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[5\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold326 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[40\] vssd1 vssd1
+ vccd1 vccd1 net1740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 team_05_WB.instance_to_wrap.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 net1751
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[16\] vssd1 vssd1
+ vccd1 vccd1 net1762 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09930_ _05938_ _05958_ vssd1 vssd1 vccd1 vccd1 _05959_ sky130_fd_sc_hd__or2_1
X_17039_ clknet_leaf_136_wb_clk_i _02669_ _00735_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold359 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[42\] vssd1 vssd1
+ vccd1 vccd1 net1773 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09365__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout806 net809 vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__clkbuf_8
X_09861_ _05888_ _05889_ vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__nand2_2
Xfanout817 _04388_ vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__buf_2
Xfanout828 _04383_ vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11172__A2 _07115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout839 net840 vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__buf_4
XANTENNA__08573__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08812_ _04878_ net377 vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__and2b_2
XANTENNA__12630__S _03682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09792_ _05208_ _05236_ vssd1 vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__nand2_1
Xhold1004 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1015 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2429 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1026 net146 vssd1 vssd1 vccd1 vccd1 net2440 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09117__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1037 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2451 sky130_fd_sc_hd__dlygate4sd3_1
X_08743_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[21\]
+ net653 _04814_ vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__a21o_1
Xhold1048 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net2462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08325__B1 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08674_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[23\]
+ net769 net746 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_159_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1090_A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13461__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout446_A net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11632__B1 _07354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10386__A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout613_A _04319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09226_ _05271_ _05273_ _05275_ _05277_ vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__or4_1
XFILLER_0_134_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09157_ net1022 _04268_ vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__and2b_2
XFILLER_0_115_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout401_X net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12805__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08108_ net1028 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[7\]
+ net975 _04203_ vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09088_ _05123_ _05144_ vssd1 vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_4_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_169_Right_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout982_A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08039_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[5\] vssd1
+ vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__inv_2
XANTENNA__10325__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold860 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold871 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2296 sky130_fd_sc_hd__dlygate4sd3_1
X_11050_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[3\] net566 _07017_
+ _07018_ vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__a22o_1
Xhold893 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2307 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09356__A2 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout770_X net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08564__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout868_X net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13636__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10001_ _06028_ _06029_ vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__nand2_1
XANTENNA__12360__B2 _07474_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12540__S net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14321__A net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09108__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08316__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1560 team_05_WB.instance_to_wrap.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 net2974
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14740_ net1066 vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__inv_2
X_11952_ _07754_ _07755_ _07763_ net343 vssd1 vssd1 vccd1 vccd1 _07764_ sky130_fd_sc_hd__o31a_1
XFILLER_0_93_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10903_ _04170_ net960 vssd1 vssd1 vccd1 vccd1 _06898_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_28_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14671_ net1233 vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11883_ _07692_ _07693_ _07688_ vssd1 vssd1 vccd1 vccd1 _07695_ sky130_fd_sc_hd__or3b_2
XANTENNA__13371__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16410_ clknet_leaf_30_wb_clk_i _02040_ _00106_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13622_ net2347 _06737_ net392 vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__mux2_1
X_17390_ clknet_leaf_57_wb_clk_i net1439 _01086_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10834_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[6\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06831_ sky130_fd_sc_hd__or2_1
XFILLER_0_156_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09816__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08318__X _04400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16341_ net1118 vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__inv_2
X_13553_ net2414 net315 net402 vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10765_ net369 _06629_ _06762_ net348 vssd1 vssd1 vccd1 vccd1 _06763_ sky130_fd_sc_hd__a211o_1
XFILLER_0_125_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12504_ net1630 _03650_ net210 vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16272_ net1124 vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__inv_2
XFILLER_0_164_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13484_ net294 net2016 net411 vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__mux2_1
X_10696_ _06628_ _06697_ net529 vssd1 vssd1 vccd1 vccd1 _06698_ sky130_fd_sc_hd__mux2_1
X_18011_ clknet_leaf_83_wb_clk_i _03350_ _01707_ vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__dfrtp_1
X_15223_ net1103 vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__inv_2
X_12435_ net1699 _07836_ _03667_ vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__mux2_1
XANTENNA__12715__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15154_ net1240 vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__inv_2
XANTENNA__09595__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12366_ net1863 net500 net217 vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_136_Right_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14105_ net910 _03970_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[10\]
+ sky130_fd_sc_hd__nor2_1
X_11317_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[16\] _07106_
+ _07108_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[88\] _07268_
+ vssd1 vssd1 vccd1 vccd1 _07276_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15085_ net1081 vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12297_ _07947_ _07959_ _03553_ vssd1 vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__a21bo_1
XANTENNA_output75_A net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14036_ _03904_ _03905_ vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__nand2_1
XANTENNA__09347__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11248_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[19\] _07106_
+ _07127_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[123\] _07209_
+ vssd1 vssd1 vccd1 vccd1 _07210_ sky130_fd_sc_hd__a221o_1
XANTENNA__14340__A2 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12351__A1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[23\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13546__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12450__S net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11179_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[7\] _07092_ _07127_
+ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[127\] _07144_ vssd1
+ vssd1 vccd1 vccd1 _07145_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15987_ net1114 vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__inv_2
XANTENNA__08307__B1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17726_ clknet_leaf_87_wb_clk_i _03069_ _01422_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[36\]
+ sky130_fd_sc_hd__dfrtp_1
X_14938_ net1055 vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_79 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17657_ clknet_leaf_41_wb_clk_i _03000_ _01353_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.next_next_data_read
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_65_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16158__A net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14869_ net1059 vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__inv_2
XANTENNA__13281__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11590__A team_05_WB.instance_to_wrap.wishbone.curr_state\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16608_ clknet_leaf_132_wb_clk_i _02238_ _00304_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_08390_ _04467_ _04469_ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__or2_4
XFILLER_0_174_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17588_ clknet_leaf_73_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[25\]
+ _01284_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13603__A1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10417__B2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11614__B1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16539_ clknet_leaf_189_wb_clk_i _02169_ _00235_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18327__1318 vssd1 vssd1 vccd1 vccd1 _18327__1318/HI net1318 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_154_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11589__X _07470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09011_ _05065_ _05067_ _05069_ _05071_ vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__or4_1
X_18209_ clknet_leaf_35_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[30\]
+ _01904_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_171_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12625__S net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold101 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[10\]
+ vssd1 vssd1 vccd1 vccd1 net1515 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[7\]
+ vssd1 vssd1 vccd1 vccd1 net1526 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold123 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[27\]
+ vssd1 vssd1 vccd1 vccd1 net1537 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold134 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[21\]
+ vssd1 vssd1 vccd1 vccd1 net1548 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08794__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold145 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[19\]
+ vssd1 vssd1 vccd1 vccd1 net1559 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold156 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[5\]
+ vssd1 vssd1 vccd1 vccd1 net1570 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold167 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[31\]
+ vssd1 vssd1 vccd1 vccd1 net1581 sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ _05531_ net373 vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__nor2_1
Xhold178 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[30\]
+ vssd1 vssd1 vccd1 vccd1 net1592 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09338__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout603 net605 vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__clkbuf_8
Xhold189 net114 vssd1 vssd1 vccd1 vccd1 net1603 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout614 _04318_ vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout396_A _03731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout625 net628 vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08546__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13456__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout636 _04312_ vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__clkbuf_8
X_09844_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[20\]
+ net818 net771 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[20\]
+ _05874_ vssd1 vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__a221o_1
Xfanout647 _04310_ vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__buf_4
Xfanout658 net659 vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1103_A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11696__A3 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[18\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout669 net671 vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__clkbuf_8
X_09775_ net370 _05596_ vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__xnor2_4
XTAP_TAPCELL_ROW_126_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08726_ _04777_ _04797_ vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08657_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[23\]
+ net600 _04730_ net721 vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout351_X net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13191__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout828_A _04383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout449_X net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08588_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[25\]
+ net831 net770 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18283__A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout616_X net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10550_ net513 _06133_ _06146_ _06559_ vssd1 vssd1 vccd1 vccd1 _06560_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_63_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09209_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[10\]
+ net836 net822 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12535__S net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10481_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[15\] _06093_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06495_ sky130_fd_sc_hd__a21oi_1
XANTENNA__14316__A net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12220_ _08021_ _03514_ _08010_ vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12151_ _07915_ _07916_ _07918_ _07960_ _07961_ vssd1 vssd1 vccd1 vccd1 _07963_ sky130_fd_sc_hd__a2111o_1
X_11102_ _07038_ _07059_ _07068_ _07031_ vssd1 vssd1 vccd1 vccd1 _07069_ sky130_fd_sc_hd__a31o_1
XFILLER_0_124_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_5__f_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12082_ net547 _07522_ vssd1 vssd1 vccd1 vccd1 _07894_ sky130_fd_sc_hd__nand2_2
Xhold690 team_05_WB.instance_to_wrap.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 net2104
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08537__B1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13366__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15910_ net1268 vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__inv_2
X_11033_ _07004_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[6\] net569
+ vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__mux2_1
XANTENNA__09734__C1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16890_ clknet_leaf_11_wb_clk_i _02520_ _00586_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15841_ net1270 vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_138_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_138_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_86_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15772_ net1299 vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__inv_2
X_12984_ net289 net2712 net464 vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__mux2_1
Xhold1390 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2804 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_26_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09501__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17511_ clknet_leaf_113_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[14\]
+ _01207_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[14\]
+ sky130_fd_sc_hd__dfrtp_2
X_11935_ _07687_ _07746_ _07710_ net343 vssd1 vssd1 vccd1 vccd1 _07747_ sky130_fd_sc_hd__o211a_1
X_14723_ net1197 vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__inv_2
XANTENNA__09799__B _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17442_ clknet_leaf_65_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[10\]
+ _01138_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_14654_ net1054 vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__inv_2
X_11866_ _07650_ _07677_ vssd1 vssd1 vccd1 vccd1 _07678_ sky130_fd_sc_hd__nand2_2
XFILLER_0_39_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13605_ net2040 net257 net392 vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__mux2_1
X_10817_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[13\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06814_ sky130_fd_sc_hd__or2_1
X_17373_ clknet_leaf_79_wb_clk_i net1419 _01069_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08068__A2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[27\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14585_ net1051 vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_60_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11797_ _07608_ _07588_ _07585_ vssd1 vssd1 vccd1 vccd1 _07609_ sky130_fd_sc_hd__mux2_2
XFILLER_0_171_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16324_ net1139 vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__inv_2
X_13536_ net2754 net226 net401 vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__mux2_1
X_10748_ net512 _06006_ _06014_ _06746_ vssd1 vssd1 vccd1 vccd1 _06747_ sky130_fd_sc_hd__a31o_1
XFILLER_0_152_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16255_ net1138 vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12445__S _03670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13467_ net238 net2184 net410 vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10679_ _05509_ net510 net333 _06207_ _06677_ vssd1 vssd1 vccd1 vccd1 _06682_ sky130_fd_sc_hd__o221a_1
XFILLER_0_129_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15206_ net1209 vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__inv_2
X_12418_ _03620_ net1758 _03668_ vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16186_ net1134 vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13398_ net2042 net218 net419 vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12572__A1 _07816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08776__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15137_ net1228 vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__inv_2
X_12349_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[20\] net996 _03616_
+ vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__a21o_4
XFILLER_0_11_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Left_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15068_ net1083 vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12324__A1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[19\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13276__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08528__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14019_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[7\] _03843_ _03888_
+ vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_leaf_65_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10335__B1 _06355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09560_ net369 _05596_ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_104_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08511_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[27\]
+ net830 net757 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17709_ clknet_leaf_91_wb_clk_i _03052_ _01405_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[83\]
+ sky130_fd_sc_hd__dfrtp_1
X_09491_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[4\]
+ net592 _05526_ _05530_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[4\]
+ sky130_fd_sc_hd__o22a_4
XFILLER_0_77_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11524__S net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08700__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08442_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[28\]
+ net670 net613 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[28\]
+ _04520_ vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_121_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09256__A1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[27\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08373_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[30\]
+ net827 net746 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_173_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1053_A net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout409_A _03728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09559__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12563__A1 _03663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_52_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1220_A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14304__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[31\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout680_A _04301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout400 net401 vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12315__A1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[21\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08519__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout411 _03728_ vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__buf_4
XANTENNA__13186__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout778_A net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout422 net423 vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__buf_6
XANTENNA_fanout399_X net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout433 _03722_ vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__clkbuf_4
Xfanout444 net447 vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__buf_6
Xfanout455 _03713_ vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__buf_4
XANTENNA__09192__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout466 _03710_ vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__buf_6
Xfanout477 net479 vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__buf_6
X_09827_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[20\]
+ net594 _05857_ net719 vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__a211o_1
XANTENNA__09731__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout488 _03700_ vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__buf_6
Xfanout499 _03696_ vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08300__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09758_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[0\]
+ net880 net873 net868 vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__and4_1
XFILLER_0_154_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08709_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[22\]
+ net796 net746 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[22\]
+ _04781_ vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_61_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout733_X net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09689_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[1\]
+ net625 _05706_ _05711_ _05712_ vssd1 vssd1 vccd1 vccd1 _05722_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10839__A team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11434__S net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11720_ _07519_ _07525_ vssd1 vssd1 vccd1 vccd1 _07532_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_81_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout900_X net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11651_ net11 net991 net918 net2954 vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__a22o_1
XFILLER_0_166_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10602_ _05816_ _05820_ vssd1 vssd1 vccd1 vccd1 _06609_ sky130_fd_sc_hd__xnor2_2
X_14370_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[13\] _04272_
+ net554 vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__a21o_1
X_11582_ net2051 net1005 _07371_ net357 vssd1 vssd1 vccd1 vccd1 _03331_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13321_ net2439 net320 net429 vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10533_ _06504_ _06543_ net518 vssd1 vssd1 vccd1 vccd1 _06544_ sky130_fd_sc_hd__mux2_1
XANTENNA__08470__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_70_Left_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16040_ net1284 vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__inv_2
X_13252_ net298 net2478 net439 vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__mux2_1
XANTENNA_input74_A wbs_we_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10464_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[17\] net904 _06475_
+ _06478_ vssd1 vssd1 vccd1 vccd1 _06479_ sky130_fd_sc_hd__a211o_1
X_12203_ net547 _07735_ vssd1 vssd1 vccd1 vccd1 _08015_ sky130_fd_sc_hd__nand2_2
X_13183_ net299 net2181 net443 vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__mux2_1
X_10395_ _06237_ _06412_ net370 vssd1 vssd1 vccd1 vccd1 _06413_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12134_ _07893_ _07898_ _07900_ _07944_ _07945_ vssd1 vssd1 vccd1 vccd1 _07946_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_20_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17991_ clknet_leaf_83_wb_clk_i _03330_ _01687_ vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13096__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12065_ _07478_ _07870_ _07872_ _07875_ _07868_ vssd1 vssd1 vccd1 vccd1 _07877_ sky130_fd_sc_hd__a41o_1
X_16942_ clknet_leaf_177_wb_clk_i _02572_ _00638_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10317__B1 _06338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18326__1317 vssd1 vssd1 vccd1 vccd1 _18326__1317/HI net1317 sky130_fd_sc_hd__conb_1
X_11016_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[9\] net569 _06990_
+ vssd1 vssd1 vccd1 vccd1 _03415_ sky130_fd_sc_hd__a21o_1
X_16873_ clknet_leaf_20_wb_clk_i _02503_ _00569_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08210__C net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08930__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15824_ net1272 vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_149_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15755_ net1304 vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__inv_2
X_12967_ net225 net2472 net466 vssd1 vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14706_ net1232 vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__inv_2
X_11918_ _07729_ _07695_ _07689_ vssd1 vssd1 vccd1 vccd1 _07730_ sky130_fd_sc_hd__mux2_2
X_15686_ net1157 vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12898_ net219 net2955 net475 vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17425_ clknet_leaf_65_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[25\]
+ _01121_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14637_ net1084 vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__inv_2
X_11849_ _07660_ vssd1 vssd1 vccd1 vccd1 _07661_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15340__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17356_ clknet_leaf_34_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[20\]
+ _01052_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_14568_ net1223 vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_35_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12683__B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11596__A2 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_109_Left_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16307_ net1164 vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__inv_2
X_13519_ net2383 net319 net405 vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__mux2_1
XANTENNA__12028__X _07840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17287_ clknet_leaf_199_wb_clk_i _02917_ _00983_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_14499_ net1207 vssd1 vssd1 vccd1 vccd1 _00129_ sky130_fd_sc_hd__inv_2
XANTENNA__08461__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload10 clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload10/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload21 clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload21/Y sky130_fd_sc_hd__inv_6
X_16238_ net1135 vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload32 clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload32/Y sky130_fd_sc_hd__clkinv_8
Xclkload43 clknet_leaf_192_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload43/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_113_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08749__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload54 clknet_leaf_177_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload54/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_3_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload65 clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload65/Y sky130_fd_sc_hd__inv_16
Xclkload76 clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload76/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_77_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16169_ net1143 vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__inv_2
Xclkload87 clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload87/Y sky130_fd_sc_hd__inv_4
XANTENNA__12903__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08213__A2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload98 clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload98/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_149_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08991_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[15\]
+ net841 _05052_ net853 vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__a211o_1
XANTENNA_clkbuf_leaf_188_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11519__S net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10308__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_118_Left_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09174__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire534_X net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_4__f_wb_clk_i_X clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09612_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[2\]
+ net880 net875 net870 vssd1 vssd1 vccd1 vccd1 _05647_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_3_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09543_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[3\]
+ net691 net624 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout261_A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17503__Q team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12577__C _07840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09474_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[4\]
+ net823 net757 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[4\]
+ _05513_ vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08425_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[29\]
+ net842 net805 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[29\]
+ _04492_ vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09229__A1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1170_A net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08356_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[30\]
+ net708 net661 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload4 clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload4/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_73_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08988__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08287_ _04236_ _04240_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[23\]
+ _04149_ _04230_ vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_33_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08452__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1056_X net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout895_A net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12813__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08204__A2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10180_ _06205_ _06206_ net526 vssd1 vssd1 vccd1 vccd1 _06207_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout683_X net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1206 net1211 vssd1 vssd1 vccd1 vccd1 net1206 sky130_fd_sc_hd__buf_2
Xfanout1217 net1220 vssd1 vssd1 vccd1 vccd1 net1217 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout230 _06367_ vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__clkbuf_2
Xfanout1228 net1234 vssd1 vssd1 vccd1 vccd1 net1228 sky130_fd_sc_hd__buf_4
Xfanout241 _06318_ vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08311__B net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09165__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1239 net1240 vssd1 vssd1 vccd1 vccd1 net1239 sky130_fd_sc_hd__clkbuf_4
Xfanout252 net253 vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_31_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout263 net266 vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__buf_2
XANTENNA_fanout850_X net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout274 net277 vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__clkbuf_2
Xfanout285 _06555_ vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout948_X net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08912__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13644__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout296 net297 vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__clkbuf_2
X_13870_ net1583 net983 _03771_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[6\]
+ sky130_fd_sc_hd__o21a_1
X_12821_ net317 net2720 net485 vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__mux2_1
XANTENNA__11672__B net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15540_ net1133 vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__inv_2
XANTENNA__10078__A2 _06106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12752_ net303 net2332 net494 vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11703_ net548 _07507_ _07514_ vssd1 vssd1 vccd1 vccd1 _07515_ sky130_fd_sc_hd__or3_1
XFILLER_0_96_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15471_ net1166 vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__inv_2
X_12683_ net2953 net339 vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__and2_1
XANTENNA__08691__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14422_ net1101 vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__inv_2
X_17210_ clknet_leaf_13_wb_clk_i _02840_ _00906_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15160__A net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11634_ team_05_WB.instance_to_wrap.wishbone.curr_state\[1\] net1 vssd1 vssd1 vccd1
+ vccd1 _07481_ sky130_fd_sc_hd__and2_1
X_18319__1411 vssd1 vssd1 vccd1 vccd1 net1411 _18319__1411/LO sky130_fd_sc_hd__conb_1
X_18190_ clknet_leaf_40_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[11\]
+ _01885_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08979__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17141_ clknet_leaf_117_wb_clk_i _02771_ _00837_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14353_ _04072_ _04076_ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__nor2_1
X_11565_ net920 _07354_ _07425_ net1007 net1584 vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__a32o_1
XANTENNA__08443__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13304_ net2145 net231 net429 vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__mux2_1
X_10516_ _05103_ _06527_ vssd1 vssd1 vccd1 vccd1 _06528_ sky130_fd_sc_hd__nor2_1
X_17072_ clknet_leaf_137_wb_clk_i _02702_ _00768_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_98_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14284_ _06481_ _06500_ _06521_ _04057_ vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__and4_1
X_11496_ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[17\] _07406_ net1003
+ vssd1 vssd1 vccd1 vccd1 _07407_ sky130_fd_sc_hd__mux2_2
XFILLER_0_12_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08205__C net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13235_ net244 net2683 net439 vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__mux2_1
X_16023_ net1284 vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__inv_2
X_10447_ net2744 net265 net539 vssd1 vssd1 vccd1 vccd1 _03456_ sky130_fd_sc_hd__mux2_1
XANTENNA__10538__B1 _04275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12723__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09157__X _05212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13166_ net245 net2122 net443 vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__mux2_1
XANTENNA__11847__B _07657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10378_ _06307_ _06396_ net532 vssd1 vssd1 vccd1 vccd1 _06397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10553__A3 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12117_ _07928_ _07916_ _07915_ vssd1 vssd1 vccd1 vccd1 _07929_ sky130_fd_sc_hd__mux2_2
Xclkbuf_leaf_153_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_153_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_20_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_72_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13097_ net189 net2123 net449 vssd1 vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__mux2_1
X_17974_ clknet_leaf_108_wb_clk_i _03313_ _01670_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08221__B net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12048_ _07859_ vssd1 vssd1 vccd1 vccd1 _07860_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_144_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16925_ clknet_leaf_109_wb_clk_i _02555_ _00621_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13554__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16856_ clknet_leaf_31_wb_clk_i _02486_ _00552_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12678__B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15807_ net1294 vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__inv_2
X_16787_ clknet_leaf_167_wb_clk_i _02417_ _00483_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13999_ _03868_ _03869_ vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15738_ net1288 vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15669_ net1256 vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__inv_2
XANTENNA__10766__X _06764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08682__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[23\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15070__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08210_ net878 net871 net867 vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__and3_4
X_17408_ clknet_leaf_64_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[8\]
+ _01104_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09190_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[10\]
+ net695 net640 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__a22o_1
X_18388_ net915 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08236__X _04319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08141_ _04221_ _04225_ _04226_ vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__and3b_1
XFILLER_0_71_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17339_ clknet_leaf_42_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[3\]
+ _01035_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08072_ net1024 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[25\]
+ net969 _04185_ vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__a22o_1
Xclkload110 clknet_leaf_162_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload110/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload121 clknet_leaf_167_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload121/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_116_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload132 clknet_leaf_142_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload132/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__12518__A1 _03646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload143 clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload143/Y sky130_fd_sc_hd__clkinv_2
Xclkload154 clknet_leaf_72_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload154/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload165 clknet_leaf_82_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload165/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_168_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12633__S net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload176 clknet_leaf_108_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload176/X sky130_fd_sc_hd__clkbuf_4
Xclkload187 clknet_leaf_96_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload187/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_168_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09395__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_126_Left_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08974_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[27\] net967
+ net955 _05036_ _04345_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[15\]
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1016_A _04347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold16 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[29\]
+ vssd1 vssd1 vccd1 vccd1 net1430 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold27 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[14\]
+ vssd1 vssd1 vccd1 vccd1 net1441 sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[13\] vssd1 vssd1
+ vccd1 vccd1 net1452 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[8\]
+ vssd1 vssd1 vccd1 vccd1 net1463 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13464__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout476_A net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09526_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[3\]
+ net752 net741 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_135_Left_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09457_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[5\]
+ net839 net835 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[5\]
+ _05491_ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout431_X net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout810_A net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09870__A1 _05888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12808__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08673__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout908_A net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11009__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08408_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[29\]
+ net676 net628 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[29\]
+ _04475_ vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09388_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[6\]
+ net699 net673 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[6\]
+ _05424_ vssd1 vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__a221o_1
XFILLER_0_136_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08339_ net950 net934 net931 vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__and3_4
X_18325__1316 vssd1 vssd1 vccd1 vccd1 _18325__1316/HI net1316 sky130_fd_sc_hd__conb_1
XFILLER_0_74_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08425__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11350_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[7\] net508 net359
+ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[3\] vssd1 vssd1 vccd1
+ vccd1 _03390_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10301_ net890 _05988_ _06322_ _06321_ vssd1 vssd1 vccd1 vccd1 _06323_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout898_X net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13639__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11281_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[114\] _07104_
+ _07111_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[106\] vssd1
+ vssd1 vccd1 vccd1 _07242_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13020_ net304 net2248 net462 vssd1 vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__mux2_1
XANTENNA__09386__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10232_ _06255_ _06256_ net372 vssd1 vssd1 vccd1 vccd1 _06257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11193__B1 _07127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_1_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1003 _07345_ vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__clkbuf_4
X_10163_ _06069_ _06076_ net514 vssd1 vssd1 vccd1 vccd1 _06190_ sky130_fd_sc_hd__mux2_1
Xfanout1014 _04371_ vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__clkbuf_4
Xfanout1025 net1026 vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__buf_2
XANTENNA__09138__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1036 team_05_WB.instance_to_wrap.total_design.core.disable_pc vssd1 vssd1 vccd1
+ vccd1 net1036 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_50_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input37_A gpio_in[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1047 team_05_WB.instance_to_wrap.total_design.core.program_count.ALU_out_reg
+ vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__buf_2
X_14971_ net1095 vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__inv_2
X_10094_ _06120_ _06121_ vssd1 vssd1 vccd1 vccd1 _06122_ sky130_fd_sc_hd__or2_1
Xfanout1058 net1064 vssd1 vssd1 vccd1 vccd1 net1058 sky130_fd_sc_hd__buf_4
XANTENNA__13374__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1069 net1108 vssd1 vssd1 vccd1 vccd1 net1069 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16710_ clknet_leaf_116_wb_clk_i _02340_ _00406_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13922_ team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.next_next_data_read
+ _03684_ vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__nand2_2
X_17690_ clknet_leaf_94_wb_clk_i _03033_ _01386_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[64\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16641_ clknet_leaf_149_wb_clk_i _02271_ _00337_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13853_ net1459 net582 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[31\]
+ sky130_fd_sc_hd__and2_1
X_12804_ net232 net2961 net487 vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16572_ clknet_leaf_157_wb_clk_i _02202_ _00268_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13784_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[13\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[12\] team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[15\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[14\] vssd1
+ vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__or4_1
X_10996_ _06819_ _06859_ _06818_ vssd1 vssd1 vccd1 vccd1 _06974_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_69_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18311_ net1403 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
XANTENNA__09310__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15523_ net1171 vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__inv_2
XANTENNA__10456__C1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12735_ net234 net2437 net494 vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__mux2_1
XANTENNA__12718__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08664__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18242_ clknet_leaf_68_wb_clk_i net1522 _01937_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15454_ net1156 vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__inv_2
X_12666_ net2946 net341 vssd1 vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09600__B net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13945__B1 _07451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14405_ net1503 vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__clkbuf_1
X_11617_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[12\] net999 vssd1
+ vssd1 vccd1 vccd1 _07479_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18173_ clknet_leaf_45_wb_clk_i _03472_ _01868_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.key_counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_137_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12597_ net1830 _03663_ _03680_ vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_137_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15385_ net1058 vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__inv_2
XANTENNA__08416__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10759__B1 _06051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08216__B net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17124_ clknet_leaf_183_wb_clk_i _02754_ _00820_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11548_ _07407_ _07392_ _07394_ _07441_ vssd1 vssd1 vccd1 vccd1 _07459_ sky130_fd_sc_hd__and4b_1
X_14336_ net349 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[9\]
+ _05351_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[8\] vssd1
+ vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_135_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold508 net85 vssd1 vssd1 vccd1 vccd1 net1922 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13549__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14267_ team_05_WB.instance_to_wrap.total_design.keypad0.counter\[0\] team_05_WB.instance_to_wrap.total_design.keypad0.counter\[1\]
+ team_05_WB.instance_to_wrap.total_design.keypad0.counter\[2\] vssd1 vssd1 vccd1
+ vccd1 _04047_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12453__S net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17055_ clknet_leaf_156_wb_clk_i _02685_ _00751_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold519 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[7\]
+ vssd1 vssd1 vccd1 vccd1 net1933 sky130_fd_sc_hd__dlygate4sd3_1
X_11479_ _07367_ _07389_ _07368_ _07363_ _07374_ vssd1 vssd1 vccd1 vccd1 _07390_ sky130_fd_sc_hd__o2111ai_4
XFILLER_0_111_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18299__1391 vssd1 vssd1 vccd1 vccd1 net1391 _18299__1391/LO sky130_fd_sc_hd__conb_1
X_16006_ net1112 vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__inv_2
X_13218_ _06637_ net353 _03718_ vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__o21ai_1
XANTENNA__14370__B1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14198_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[6\] _04000_
+ vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11184__B1 _07108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ net286 net2945 net444 vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1208 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2622 sky130_fd_sc_hd__dlygate4sd3_1
X_17957_ clknet_leaf_107_wb_clk_i _03296_ _01653_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__dfrtp_1
Xhold1219 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2633 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13284__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16908_ clknet_leaf_7_wb_clk_i _02538_ _00604_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08690_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[22\]
+ net708 net637 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[22\]
+ _04761_ vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__a221o_1
X_17888_ clknet_leaf_104_wb_clk_i _03231_ _01584_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16839_ clknet_leaf_202_wb_clk_i _02469_ _00535_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12436__A0 _03641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_50_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09311_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[8\]
+ net762 net747 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__a22o_1
XANTENNA__12628__S net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11532__S net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09242_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[9\]
+ net693 net623 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[9\]
+ _05290_ vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_157_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10656__B net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09173_ _05221_ _05223_ _05225_ _05226_ vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__or4_2
XANTENNA__08407__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08124_ net154 net153 vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09080__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13459__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08055_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[11\] vssd1 vssd1
+ vccd1 vccd1 _04175_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1133_A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout593_A _04368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1300_A net1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1019_X net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18318__1410 vssd1 vssd1 vccd1 vccd1 net1410 _18318__1410/LO sky130_fd_sc_hd__conb_1
X_08957_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[15\]
+ net676 net652 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout760_A net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13194__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout858_A net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout479_X net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08888_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[17\]
+ net806 net745 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__a22o_1
XANTENNA__09540__B1 _05556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10150__A1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout646_X net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11008__A _04170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10850_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[3\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[3\]
+ _06846_ vssd1 vssd1 vccd1 vccd1 _06847_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09509_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[4\]
+ net661 _05547_ net721 vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__a211o_1
XFILLER_0_6_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12538__S net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10781_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[29\] net1040 vssd1
+ vssd1 vccd1 vccd1 _06778_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout813_X net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08646__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12520_ net1653 _03610_ net209 vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12451_ net1733 _03610_ net213 vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11402_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[16\] _07330_
+ vssd1 vssd1 vccd1 vccd1 _07332_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15170_ net1204 vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__inv_2
X_12382_ net1755 _03612_ net216 vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09071__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14121_ _03983_ _03984_ vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13369__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11333_ _07288_ _07290_ vssd1 vssd1 vccd1 vccd1 _07291_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_10_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09359__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14052_ _03890_ _03898_ _03920_ vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_132_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11264_ _07219_ _07221_ _07223_ _07225_ vssd1 vssd1 vccd1 vccd1 _07226_ sky130_fd_sc_hd__or4_1
XFILLER_0_123_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11166__B1 _07128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13003_ net236 net2688 net462 vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10215_ _06003_ _06229_ _06240_ net338 vssd1 vssd1 vccd1 vccd1 _06241_ sky130_fd_sc_hd__o22a_1
X_11195_ _07156_ _07158_ _07159_ vssd1 vssd1 vccd1 vccd1 _07160_ sky130_fd_sc_hd__or3_1
XFILLER_0_24_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17811_ clknet_leaf_74_wb_clk_i _03154_ _01507_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10146_ _04573_ net363 vssd1 vssd1 vccd1 vccd1 _06174_ sky130_fd_sc_hd__nand2_1
X_17742_ clknet_leaf_87_wb_clk_i _03085_ _01438_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[52\]
+ sky130_fd_sc_hd__dfrtp_1
X_10077_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[31\] net904 net968
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[31\] _06105_ vssd1
+ vssd1 vccd1 vccd1 _06106_ sky130_fd_sc_hd__a221o_2
X_14954_ net1113 vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_89_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13905_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[24\]
+ net559 net575 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[24\]
+ net986 vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__a221o_1
XFILLER_0_89_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17673_ clknet_leaf_100_wb_clk_i _03016_ _01369_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[111\]
+ sky130_fd_sc_hd__dfrtp_1
X_14885_ net1196 vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__inv_2
XANTENNA__08885__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload2_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16624_ clknet_leaf_124_wb_clk_i _02254_ _00320_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13836_ net1486 net578 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[14\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_43_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13091__A0 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16555_ clknet_leaf_186_wb_clk_i _02185_ _00251_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13767_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[25\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[24\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[27\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[26\]
+ vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__or4_1
XANTENNA__12448__S _03670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10979_ _06960_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[16\] net564
+ vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__mux2_1
XANTENNA__08637__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11205__X _07169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15506_ net1173 vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__inv_2
X_12718_ net320 net2685 net497 vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_63_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16486_ clknet_leaf_116_wb_clk_i _02116_ _00182_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13698_ team_05_WB.instance_to_wrap.wishbone.curr_state\[1\] _04169_ _07490_ team_05_WB.instance_to_wrap.wishbone.curr_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18225_ clknet_leaf_66_wb_clk_i net1481 _01920_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_135_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15437_ net1164 vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__inv_2
X_12649_ team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.next_next_data_read
+ _03687_ _03685_ vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__o21a_1
XFILLER_0_109_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09598__B1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18156_ clknet_leaf_160_wb_clk_i _03459_ _01852_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_15368_ net1218 vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08514__X team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[27\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09062__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13279__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17107_ clknet_leaf_166_wb_clk_i _02737_ _00803_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold305 net122 vssd1 vssd1 vccd1 vccd1 net1719 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14319_ _04818_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[21\]
+ net360 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[20\] _04091_
+ vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__a221o_1
Xhold316 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[69\] vssd1 vssd1
+ vccd1 vccd1 net1730 sky130_fd_sc_hd__dlygate4sd3_1
X_18087_ clknet_leaf_79_wb_clk_i _03410_ _01783_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15299_ net1206 vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__inv_2
Xhold327 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[68\] vssd1 vssd1
+ vccd1 vccd1 net1741 sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[45\] vssd1 vssd1
+ vccd1 vccd1 net1752 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold349 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[16\] vssd1 vssd1
+ vccd1 vccd1 net1763 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17038_ clknet_leaf_173_wb_clk_i _02668_ _00734_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09860_ _04839_ _05881_ _05885_ vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__a21boi_2
Xfanout807 net809 vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12911__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout818 net821 vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_110_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout829 net832 vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__clkbuf_8
X_08811_ _04879_ vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__inv_2
XANTENNA__09770__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09791_ _05284_ _05821_ _05282_ vssd1 vssd1 vccd1 vccd1 _05822_ sky130_fd_sc_hd__a21o_1
XANTENNA__10380__A1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10380__B2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1005 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 net2419 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11527__S net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1016 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 net2430 sky130_fd_sc_hd__dlygate4sd3_1
X_08742_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[21\]
+ net622 net618 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[21\]
+ net719 vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__a221o_1
XANTENNA__09064__Y _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1027 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net2441 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1038 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2452 sky130_fd_sc_hd__dlygate4sd3_1
X_18324__1315 vssd1 vssd1 vccd1 vccd1 _18324__1315/HI net1315 sky130_fd_sc_hd__conb_1
Xhold1049 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2463 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09522__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08673_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[23\]
+ net819 net807 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[23\]
+ _04746_ vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__a221o_1
XFILLER_0_139_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12409__A0 _03651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08628__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout341_A _03693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17511__Q team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[14\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1083_A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout439_A _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11632__A1 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10386__B _06404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09225_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[10\]
+ net849 _05276_ net853 vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__a211o_1
XFILLER_0_57_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout606_A _04320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09156_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[7\] net1022
+ _04268_ net966 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__a32o_1
XANTENNA__09053__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08107_ net1028 net2771 vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__and2b_1
XANTENNA__13189__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09087_ net572 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[13\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[13\] vssd1 vssd1 vccd1
+ vccd1 _05144_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08800__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08038_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[12\] vssd1 vssd1
+ vccd1 vccd1 _04160_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold850 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2264 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout975_A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold861 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net2275 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout596_X net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold872 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net2286 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11699__A1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[20\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold883 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2297 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12821__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold894 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 net2308 sky130_fd_sc_hd__dlygate4sd3_1
X_10000_ _05165_ net362 vssd1 vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__nand2_1
XANTENNA__10371__A1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout763_X net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14321__B team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[23\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09989_ _05208_ net361 vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__or2_1
XFILLER_0_157_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1550 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 net2964 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1561 team_05_WB.instance_to_wrap.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 net2975
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11951_ _07753_ _07760_ vssd1 vssd1 vccd1 vccd1 _07763_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout930_X net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11320__B1 _07105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08867__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13652__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10902_ _06777_ _06778_ vssd1 vssd1 vccd1 vccd1 _06897_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_28_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14670_ net1187 vssd1 vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__inv_2
X_11882_ _07659_ _07663_ vssd1 vssd1 vccd1 vccd1 _07694_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18298__1390 vssd1 vssd1 vccd1 vccd1 net1390 _18298__1390/LO sky130_fd_sc_hd__conb_1
XFILLER_0_79_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10833_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[6\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06830_ sky130_fd_sc_hd__nand2_1
X_13621_ net2565 net310 net392 vssd1 vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08619__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16340_ net1124 vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13552_ net2465 net317 net401 vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__mux2_1
X_10764_ net526 _06697_ _06761_ net370 vssd1 vssd1 vccd1 vccd1 _06762_ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09292__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12503_ net1849 _07816_ _03673_ vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__mux2_1
X_16271_ net1113 vssd1 vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__inv_2
X_13483_ net301 net2381 net411 vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10695_ _06661_ _06696_ net516 vssd1 vssd1 vccd1 vccd1 _06697_ sky130_fd_sc_hd__mux2_1
X_18010_ clknet_leaf_64_wb_clk_i _03349_ _01706_ vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__dfrtp_1
XANTENNA__13376__A1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12434_ _03650_ net1819 _03668_ vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__mux2_1
X_15222_ net1091 vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10583__Y _06591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13099__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12365_ _07858_ _07859_ _07863_ _03659_ vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__and4_4
XFILLER_0_152_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15153_ net1192 vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_130_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08053__Y _04173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11316_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[120\] _07099_
+ _07274_ vssd1 vssd1 vccd1 vccd1 _07275_ sky130_fd_sc_hd__a21o_1
X_14104_ net1642 net506 _03969_ vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_121_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15084_ net1071 vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__inv_2
X_12296_ _03590_ vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14035_ _03872_ _03903_ _03873_ vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__or3b_1
X_11247_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[107\] _07102_
+ _07104_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[115\] vssd1
+ vssd1 vccd1 vccd1 _07209_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_55_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09201__C1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12731__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11178_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[47\] _07091_
+ _07103_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[119\] vssd1
+ vssd1 vccd1 vccd1 _07144_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_1064 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10129_ net380 net368 vssd1 vssd1 vccd1 vccd1 _06157_ sky130_fd_sc_hd__nand2_1
X_15986_ net1128 vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_69_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09504__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17725_ clknet_leaf_101_wb_clk_i _03068_ _01421_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14937_ net1053 vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__inv_2
XANTENNA__11311__B1 _07120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13562__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17656_ clknet_leaf_39_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[23\]
+ _01352_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14868_ net1075 vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__inv_2
XANTENNA__12686__B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10758__Y _06756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11590__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16607_ clknet_leaf_155_wb_clk_i _02237_ _00303_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13819_ net1592 net969 net723 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[30\]
+ sky130_fd_sc_hd__and3_1
X_17587_ clknet_leaf_113_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[24\]
+ _01283_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14799_ net1286 vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__inv_2
X_16538_ clknet_leaf_31_wb_clk_i _02168_ _00234_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11614__A1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[14\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09283__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08491__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12906__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16469_ clknet_leaf_173_wb_clk_i _02099_ _00165_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16174__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09010_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[14\]
+ net627 net609 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[14\]
+ _05070_ vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__a221o_1
X_18208_ clknet_leaf_37_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[29\]
+ _01903_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_171_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_94_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09035__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18139_ clknet_leaf_165_wb_clk_i _03442_ _01835_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08243__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10426__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold102 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[5\]
+ vssd1 vssd1 vccd1 vccd1 net1516 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11709__C_N team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold113 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[29\]
+ vssd1 vssd1 vccd1 vccd1 net1527 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[20\]
+ vssd1 vssd1 vccd1 vccd1 net1538 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold135 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[11\]
+ vssd1 vssd1 vccd1 vccd1 net1549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[12\]
+ vssd1 vssd1 vccd1 vccd1 net1560 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold157 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[4\]
+ vssd1 vssd1 vccd1 vccd1 net1571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 net87 vssd1 vssd1 vccd1 vccd1 net1582 sky130_fd_sc_hd__dlygate4sd3_1
X_09912_ net374 _05505_ vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__and2b_1
Xhold179 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[16\]
+ vssd1 vssd1 vccd1 vccd1 net1593 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12641__S net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout604 net605 vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__clkbuf_4
Xfanout615 _04318_ vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__clkbuf_8
Xfanout626 net628 vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09843_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[20\]
+ net778 net768 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__a22o_1
Xfanout637 _04312_ vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout648 net651 vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__buf_6
Xfanout659 _04307_ vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__buf_4
XFILLER_0_77_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout389_A _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09774_ net370 _05596_ vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__nand2_1
X_08725_ _04344_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[22\]
+ _04362_ vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11302__B1 _07092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_201_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08849__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13472__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1298_A net1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08656_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[23\]
+ net688 net653 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08587_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[25\]
+ net828 net804 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[25\]
+ _04662_ vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout723_A net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1086_X net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11605__B2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[20\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10684__X _06687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08482__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout511_X net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12816__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout609_X net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09208_ _05260_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[10\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_91_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10480_ _06488_ _06493_ net538 vssd1 vssd1 vccd1 vccd1 _06494_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09026__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14316__B team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[19\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09139_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[11\]
+ net629 net602 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08314__B net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12150_ _07960_ _07961_ vssd1 vssd1 vccd1 vccd1 _07962_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10592__A1 _06049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11101_ _07063_ _07067_ vssd1 vssd1 vccd1 vccd1 _07068_ sky130_fd_sc_hd__and2_2
XANTENNA__13647__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12551__S net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12081_ _07885_ _07890_ _07892_ _07883_ vssd1 vssd1 vccd1 vccd1 _07893_ sky130_fd_sc_hd__o22ai_2
XANTENNA__12404__X _03667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold680 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net2094 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14332__A net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold691 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 net2105 sky130_fd_sc_hd__dlygate4sd3_1
X_11032_ net964 _06658_ _07003_ vssd1 vssd1 vccd1 vccd1 _07004_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13530__A1 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08330__A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15840_ net1276 vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__inv_2
XANTENNA__10895__A2 _05921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_139_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11962__Y _07774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13294__A0 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15771_ net1305 vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12983_ net291 net2693 net464 vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__mux2_1
XANTENNA__13382__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17510_ clknet_leaf_73_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[13\]
+ _01206_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[13\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold1380 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1391 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2805 sky130_fd_sc_hd__dlygate4sd3_1
X_14722_ net1228 vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__inv_2
X_11934_ _07707_ _07708_ _07712_ vssd1 vssd1 vccd1 vccd1 _07746_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09161__A _05215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17441_ clknet_leaf_65_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[9\]
+ _01137_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_178_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_178_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_14653_ net1090 vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11865_ _07669_ _07671_ _07673_ _07674_ _07675_ vssd1 vssd1 vccd1 vccd1 _07677_ sky130_fd_sc_hd__a32o_1
XFILLER_0_129_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13604_ net2553 net254 net392 vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_107_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_107_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_17372_ clknet_leaf_81_wb_clk_i net1434 _01068_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10816_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[13\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06813_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14584_ net1200 vssd1 vssd1 vccd1 vccd1 _00214_ sky130_fd_sc_hd__inv_2
X_11796_ _07582_ _07588_ vssd1 vssd1 vccd1 vccd1 _07608_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16323_ net1139 vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__inv_2
XFILLER_0_165_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13535_ net2959 net233 net402 vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10747_ net517 _06004_ _06007_ net525 vssd1 vssd1 vccd1 vccd1 _06746_ sky130_fd_sc_hd__a31o_1
XFILLER_0_83_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10280__B1 _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16254_ net1131 vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13466_ net242 net2191 net411 vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__mux2_1
XANTENNA__09017__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10678_ net524 _06612_ _06680_ vssd1 vssd1 vccd1 vccd1 _06681_ sky130_fd_sc_hd__a21o_1
X_18323__1314 vssd1 vssd1 vccd1 vccd1 _18323__1314/HI net1314 sky130_fd_sc_hd__conb_1
XFILLER_0_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15205_ net1194 vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__inv_2
X_12417_ _03644_ net1848 net214 vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__mux2_1
X_16185_ net1135 vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__inv_2
X_13397_ net2178 net189 net417 vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__mux2_1
X_15136_ net1198 vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__inv_2
X_12348_ net545 _07507_ net500 _07864_ _07914_ vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_65_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_178_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13557__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15338__A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12461__S net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12279_ _03560_ _03566_ _03570_ _03558_ vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__o22ai_2
X_15067_ net1075 vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__inv_2
XANTENNA__09725__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14018_ _03861_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[7\] vssd1
+ vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_147_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15969_ net1275 vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08510_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[27\]
+ net753 net742 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__a22o_1
XANTENNA__13292__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17708_ clknet_leaf_84_wb_clk_i _03051_ _01404_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[82\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15073__A net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09490_ _05514_ _05517_ _05528_ _05529_ vssd1 vssd1 vccd1 vccd1 _05530_ sky130_fd_sc_hd__or4_1
XFILLER_0_77_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08441_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[28\]
+ net623 net609 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__a22o_1
X_17639_ clknet_leaf_67_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[6\]
+ _01335_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_121_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08372_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[30\]
+ net816 net788 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[30\]
+ _04452_ vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__a221o_1
XFILLER_0_81_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_862 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11599__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12636__S net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08464__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09008__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout304_A _06655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1046_A net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08767__A1 _04344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13467__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12371__S net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09517__Y _05556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1213_A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13512__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout401 net403 vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__clkbuf_8
Xfanout412 _03727_ vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__buf_8
Xfanout423 _03725_ vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08150__A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout434 _03722_ vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__buf_6
XANTENNA_clkbuf_3_6_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout445 net447 vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout673_A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout456 _03712_ vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__buf_8
X_09826_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[20\]
+ net687 net598 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__a22o_1
Xfanout467 _03710_ vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__buf_4
Xfanout478 net479 vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__buf_4
Xfanout489 _03700_ vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__buf_4
XANTENNA_fanout461_X net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09757_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[0\]
+ net880 net873 net859 vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__and4_1
Xclkbuf_leaf_5_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout938_A net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08708_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[22\]
+ net839 net743 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09688_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[1\]
+ net699 _05701_ _05714_ _05716_ vssd1 vssd1 vccd1 vccd1 _05721_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09495__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09908__A_N _05165_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18067__Q net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08639_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[24\]
+ net824 net773 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[24\]
+ _04713_ vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__a221o_1
XFILLER_0_51_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout726_X net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12894__X _03706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_200_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_200_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__15711__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11650_ net12 net991 net918 net2306 vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09247__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10601_ _05820_ _05956_ _06607_ vssd1 vssd1 vccd1 vccd1 _06608_ sky130_fd_sc_hd__a21oi_1
X_11581_ net1924 net1005 _07373_ net357 vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__a22o_1
XANTENNA__11054__A2 _06729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08455__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12546__S net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13320_ net2529 net304 net429 vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__mux2_1
X_10532_ _06026_ _06028_ vssd1 vssd1 vccd1 vccd1 _06543_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10463_ net895 _06477_ _05485_ vssd1 vssd1 vccd1 vccd1 _06478_ sky130_fd_sc_hd__o21ai_1
X_13251_ net287 net2369 net436 vssd1 vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__mux2_1
XANTENNA__13200__A0 _06317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12202_ _07994_ _07997_ _08013_ _07991_ vssd1 vssd1 vccd1 vccd1 _08014_ sky130_fd_sc_hd__a22o_1
X_13182_ net286 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[10\]
+ net440 vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__mux2_1
XANTENNA_input67_A wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10394_ _06336_ _06411_ net530 vssd1 vssd1 vccd1 vccd1 _06412_ sky130_fd_sc_hd__mux2_1
XANTENNA__13377__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12133_ _07871_ _07881_ _07891_ vssd1 vssd1 vccd1 vccd1 _07945_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_36_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17990_ clknet_leaf_83_wb_clk_i _03329_ _01686_ vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12064_ _07872_ _07875_ vssd1 vssd1 vccd1 vccd1 _07876_ sky130_fd_sc_hd__nand2_1
X_16941_ clknet_leaf_158_wb_clk_i _02571_ _00637_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11015_ net963 _06609_ _06989_ vssd1 vssd1 vccd1 vccd1 _06990_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_53_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16872_ clknet_leaf_204_wb_clk_i _02502_ _00568_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08995__A _05034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout990 _07482_ vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__buf_2
X_15823_ net1290 vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_5_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15754_ net1295 vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_142_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12966_ net218 net2583 net467 vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__mux2_1
X_14705_ net1189 vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ _07695_ _07697_ vssd1 vssd1 vccd1 vccd1 _07729_ sky130_fd_sc_hd__nand2_1
X_15685_ net1156 vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__inv_2
XANTENNA__12490__A1 _03612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11293__A2 _07102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08694__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12897_ net190 net2727 net473 vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__mux2_1
XANTENNA__08219__B net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17424_ clknet_leaf_61_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[24\]
+ _01120_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14636_ net1121 vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11848_ _07656_ _07659_ vssd1 vssd1 vccd1 vccd1 _07660_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09238__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17355_ clknet_leaf_36_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[19\]
+ _01051_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08446__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12456__S net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14567_ net1242 vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__inv_2
XANTENNA__12309__X _03604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11779_ _07577_ _07578_ _07573_ vssd1 vssd1 vccd1 vccd1 _07591_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16306_ net1161 vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__inv_2
XFILLER_0_166_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13518_ net2670 net302 net405 vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__mux2_1
X_17286_ clknet_leaf_116_wb_clk_i _02916_ _00982_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14498_ net1193 vssd1 vssd1 vccd1 vccd1 _00128_ sky130_fd_sc_hd__inv_2
X_16237_ net1135 vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__inv_2
Xclkload11 clknet_leaf_195_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload11/Y sky130_fd_sc_hd__inv_6
X_13449_ net2119 net287 net412 vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__mux2_1
Xclkload22 clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload22/Y sky130_fd_sc_hd__inv_6
Xclkload33 clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload33/Y sky130_fd_sc_hd__bufinv_16
Xclkbuf_leaf_75_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload44 clknet_leaf_193_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload44/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_70_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload55 clknet_leaf_178_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload55/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16168_ net1143 vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__inv_2
Xclkload66 clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload66/Y sky130_fd_sc_hd__clkinv_8
Xclkload77 clknet_leaf_47_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload77/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__10771__Y _06768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10556__A1 _06049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09410__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload88 clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload88/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__10556__B2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload99 clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload99/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_149_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13287__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15119_ net1240 vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__inv_2
XANTENNA__10704__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16099_ net1307 vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__inv_2
X_08990_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[15\]
+ net837 net756 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_166_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10005__A net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09611_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[2\]
+ net885 net871 net857 vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_123_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09513__B net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09542_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[3\]
+ net636 net617 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09477__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11284__A2 _07110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12481__A1 _07791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09473_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[4\]
+ net807 net783 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__a22o_1
X_08424_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[29\]
+ net798 net787 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[29\]
+ _04498_ vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__a221o_1
XANTENNA__09229__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08355_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[30\]
+ net653 net603 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[30\]
+ _04434_ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12366__S net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08437__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout421_A net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1163_A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout519_A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11587__A3 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload5 clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload5/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_11_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08286_ net945 _04366_ vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__nand2_8
XFILLER_0_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13986__A _07380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout307_X net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1049_X net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout790_A net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09401__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout888_A _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13197__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1207 net1210 vssd1 vssd1 vccd1 vccd1 net1207 sky130_fd_sc_hd__buf_4
Xfanout1218 net1219 vssd1 vssd1 vccd1 vccd1 net1218 sky130_fd_sc_hd__buf_4
Xfanout220 net221 vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout676_X net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout231 _06367_ vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1229 net1234 vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__buf_2
Xfanout242 net244 vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08311__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout253 _06423_ vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__clkbuf_2
Xfanout264 net266 vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_31_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout275 net277 vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__clkbuf_2
Xfanout286 net287 vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__clkbuf_2
X_09809_ _04924_ _05839_ _04922_ vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__o21a_2
Xfanout297 _06638_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout843_X net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11445__S net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12820_ net303 net2128 net486 vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11672__C net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11275__A2 _07113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12472__A1 _03623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12751_ net296 net2708 net495 vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13660__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11702_ _07508_ _07509_ _07511_ _07513_ vssd1 vssd1 vccd1 vccd1 _07514_ sky130_fd_sc_hd__or4_1
X_15470_ net1171 vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__inv_2
X_12682_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[7\]
+ net341 vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__and2_1
XFILLER_0_166_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14421_ net1080 vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11633_ net145 net1012 _07471_ net2818 vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__a22o_1
XANTENNA__08428__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17140_ clknet_leaf_119_wb_clk_i _02770_ _00836_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14352_ _04064_ _04124_ _04075_ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__a21o_1
X_11564_ net1804 net1004 _07432_ net358 vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13303_ net2413 net236 net429 vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_98_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10515_ _04158_ _05102_ _06051_ vssd1 vssd1 vccd1 vccd1 _06527_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17071_ clknet_leaf_136_wb_clk_i _02701_ _00767_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_98_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11495_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[17\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[17\]
+ net1031 vssd1 vssd1 vccd1 vccd1 _07406_ sky130_fd_sc_hd__mux2_1
X_14283_ _06540_ _06557_ _04056_ vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_1012 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16022_ net1284 vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__inv_2
X_13234_ net224 net2687 net438 vssd1 vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__mux2_1
X_10446_ net382 _06461_ vssd1 vssd1 vccd1 vccd1 _06462_ sky130_fd_sc_hd__and2_1
XFILLER_0_150_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18260__Q team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[14\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13165_ net224 net2303 net442 vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__mux2_1
X_10377_ _06357_ _06395_ net518 vssd1 vssd1 vccd1 vccd1 _06396_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12116_ _07916_ _07918_ vssd1 vssd1 vccd1 vccd1 _07928_ sky130_fd_sc_hd__nand2_1
X_13096_ net193 net2254 net450 vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__mux2_1
X_17973_ clknet_leaf_107_wb_clk_i _03312_ _01669_ vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09156__A1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08221__C net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12047_ _07377_ _07468_ _07845_ _07369_ vssd1 vssd1 vccd1 vccd1 _07859_ sky130_fd_sc_hd__or4b_2
XTAP_TAPCELL_ROW_144_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16924_ clknet_leaf_155_wb_clk_i _02554_ _00620_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11499__C1 _07409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_193_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_193_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16855_ clknet_leaf_143_wb_clk_i _02485_ _00551_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15806_ net1297 vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_161_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_122_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_122_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16786_ clknet_leaf_127_wb_clk_i _02416_ _00482_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13998_ net978 team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[12\] vssd1
+ vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__and2_1
XANTENNA__09459__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15737_ net1267 vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12463__A1 _07797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11266__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12949_ net279 net2384 net468 vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__mux2_1
XANTENNA__08667__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13570__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10474__B1 _06333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15668_ net1256 vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17407_ clknet_leaf_65_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[7\]
+ _01103_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14619_ net1098 vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__inv_2
XANTENNA__08419__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18387_ net1369 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__buf_2
X_15599_ net1258 vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__inv_2
X_08140_ team_05_WB.instance_to_wrap.total_design.keypad0.key_counter\[2\] _04220_
+ vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17338_ clknet_leaf_36_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[2\]
+ _01034_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09092__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload100 clknet_leaf_65_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload100/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_153_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08071_ net1024 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__and2b_1
XFILLER_0_43_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload111 clknet_leaf_163_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload111/X sky130_fd_sc_hd__clkbuf_8
X_17269_ clknet_leaf_173_wb_clk_i _02899_ _00965_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12914__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload122 clknet_leaf_168_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload122/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_141_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload133 clknet_leaf_143_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload133/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload144 clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload144/Y sky130_fd_sc_hd__clkinv_2
Xclkload155 clknet_leaf_74_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload155/Y sky130_fd_sc_hd__inv_8
Xclkload166 clknet_leaf_84_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload166/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_168_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload177 clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload177/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_168_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08198__A2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload188 clknet_leaf_97_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload188/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_41_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13479__A0 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08973_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[15\] _04355_
+ vssd1 vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__xnor2_1
Xhold17 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[31\]
+ vssd1 vssd1 vccd1 vccd1 net1431 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold28 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[23\]
+ vssd1 vssd1 vccd1 vccd1 net1442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[22\] vssd1 vssd1
+ vccd1 vccd1 net1453 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1009_A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17514__Q team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[17\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout371_A net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08370__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout469_A net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09525_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[3\]
+ net793 net782 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__a22o_1
XANTENNA__11257__A2 _07096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12454__A1 _03614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08658__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1280_A net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13480__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout636_A _04312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_5_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09456_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[5\]
+ net812 net800 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[5\]
+ _05487_ vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__a221o_1
XFILLER_0_137_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11009__A2 _06603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08407_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[29\]
+ net696 net646 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[29\]
+ _04476_ vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__a221o_1
XFILLER_0_109_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09387_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[6\]
+ net669 net661 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[6\]
+ _05431_ vssd1 vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout424_X net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout803_A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10217__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08338_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[31\]
+ net746 net742 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09083__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10768__A1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09622__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08269_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[29\] _04351_
+ vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__or2_2
XFILLER_0_7_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12824__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10300_ _05898_ _05984_ _05987_ vssd1 vssd1 vccd1 vccd1 _06322_ sky130_fd_sc_hd__nor3_1
XFILLER_0_15_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11280_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[10\] _07105_
+ _07106_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[18\] _07235_
+ vssd1 vssd1 vccd1 vccd1 _07241_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout793_X net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10231_ _06046_ _06080_ net530 vssd1 vssd1 vccd1 vccd1 _06256_ sky130_fd_sc_hd__mux2_1
XANTENNA__08322__B net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10162_ _06186_ _06188_ _05924_ vssd1 vssd1 vccd1 vccd1 _06189_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_7_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1004 net1006 vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__buf_2
Xfanout1015 _04347_ vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__buf_2
XANTENNA__13655__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1026 net1036 vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_50_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1037 net1039 vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__clkbuf_2
X_14970_ net1053 vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_50_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10093_ _05596_ net366 vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__nor2_1
Xfanout1048 team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.state\[2\] vssd1
+ vssd1 vccd1 vccd1 net1048 sky130_fd_sc_hd__clkbuf_2
Xfanout1059 net1061 vssd1 vssd1 vccd1 vccd1 net1059 sky130_fd_sc_hd__buf_4
XANTENNA__09689__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13921_ team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.next_next_data_read
+ _03684_ vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__and2_1
XANTENNA__08897__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16640_ clknet_leaf_126_wb_clk_i _02270_ _00336_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13852_ net1484 net578 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[30\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_92_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10299__B _06320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12803_ net236 net2109 net486 vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__mux2_1
XANTENNA__12445__A1 _07789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11248__A2 _07106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16571_ clknet_leaf_194_wb_clk_i _02201_ _00267_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08649__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13783_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[9\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[8\] team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[11\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[10\] vssd1
+ vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__or4_1
X_10995_ net1452 net568 _06973_ vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__a21o_1
XANTENNA__09846__C1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13390__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18310_ net1402 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
X_15522_ net1170 vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12734_ net238 net2569 net495 vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18241_ clknet_leaf_59_wb_clk_i net1588 _01936_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__18255__Q team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15453_ net1147 vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__inv_2
X_12665_ net2562 net341 vssd1 vssd1 vccd1 vccd1 _02958_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08056__Y _04176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14404_ net1551 vssd1 vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__clkbuf_1
X_18172_ clknet_leaf_45_wb_clk_i _03471_ _01867_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.key_counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11616_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[12\] net997 vssd1
+ vssd1 vccd1 vccd1 _07478_ sky130_fd_sc_hd__and2_2
XFILLER_0_154_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09074__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15384_ net1244 vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__inv_2
X_12596_ net1650 _07812_ _03680_ vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10759__A1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17123_ clknet_leaf_199_wb_clk_i _02753_ _00819_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_14335_ _05256_ net534 net349 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__o2bb2a_1
X_11547_ _07453_ _07455_ _07456_ _07457_ vssd1 vssd1 vccd1 vccd1 _07458_ sky130_fd_sc_hd__or4_2
XANTENNA__08821__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12734__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold509 team_05_WB.instance_to_wrap.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 net1923
+ sky130_fd_sc_hd__dlygate4sd3_1
X_17054_ clknet_leaf_163_wb_clk_i _02684_ _00750_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_14266_ _04018_ _04046_ vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__and2_1
X_11478_ _07383_ _07387_ _07353_ vssd1 vssd1 vccd1 vccd1 _07389_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_74_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16005_ net1114 vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__inv_2
XANTENNA__14370__A1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13217_ net2521 net353 vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__nand2_1
X_10429_ _04925_ _05839_ vssd1 vssd1 vccd1 vccd1 _06445_ sky130_fd_sc_hd__xnor2_4
X_14197_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[6\] _04000_
+ vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__or2_1
XANTENNA__08232__B net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ net291 net2674 net444 vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_163_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13565__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13792__C net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13079_ net274 net2865 net455 vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__mux2_1
X_17956_ clknet_leaf_108_wb_clk_i _03295_ _01652_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__dfrtp_1
Xhold1209 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2623 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12689__B net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16907_ clknet_leaf_189_wb_clk_i _02537_ _00603_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_17887_ clknet_leaf_75_wb_clk_i _03230_ _01583_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08888__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08352__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16838_ clknet_leaf_118_wb_clk_i _02468_ _00534_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11239__A2 _07111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16769_ clknet_leaf_149_wb_clk_i _02399_ _00465_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12909__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08104__A2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15081__A net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09310_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[8\]
+ net831 net800 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09350__Y _05397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10998__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09241_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[9\]
+ net713 net697 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[9\]
+ _05291_ vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__a221o_1
XANTENNA__18392__A net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_90_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_118_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09172_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[11\]
+ net786 net764 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[11\]
+ _05216_ vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08123_ net35 net37 net36 net34 vssd1 vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__or4b_1
XFILLER_0_114_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12644__S net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout217_A _03660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08054_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[8\] vssd1 vssd1
+ vccd1 vccd1 _04174_ sky130_fd_sc_hd__inv_2
XANTENNA__17509__Q team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[12\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1126_A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13475__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13328__X _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08591__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15256__A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08956_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[15\]
+ net699 net625 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[15\]
+ _05018_ vssd1 vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__a221o_1
XANTENNA__08328__C1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08887_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[17\]
+ _04383_ net744 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[17\]
+ _04947_ vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout753_A net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09540__A1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08343__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout920_A _07352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12427__A1 _07798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12819__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout541_X net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout639_X net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09260__Y team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09508_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[4\]
+ net666 net638 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__a22o_1
XANTENNA__09701__B _05731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10780_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[29\] net1040 vssd1
+ vssd1 vccd1 vccd1 _06777_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10989__A1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09843__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09439_ _05468_ _05470_ _05480_ _05481_ vssd1 vssd1 vccd1 vccd1 _05482_ sky130_fd_sc_hd__or4_1
XANTENNA__11650__A2 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10339__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout806_X net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12450_ net1649 _03655_ net212 vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__mux2_1
XANTENNA__09056__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11401_ net1554 _07331_ vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12381_ net1701 _03614_ net216 vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__mux2_1
XANTENNA__08803__B1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14120_ _03950_ _03972_ _03982_ vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__or3b_1
X_11332_ _07286_ _07289_ vssd1 vssd1 vccd1 vccd1 _07290_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08333__A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14051_ _03918_ _03919_ vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__nor2_1
X_11263_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[19\] _07125_
+ _07130_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[99\] _07224_
+ vssd1 vssd1 vccd1 vccd1 _07225_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_91_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_45_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13002_ net240 net2118 net463 vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__mux2_1
X_10214_ _06238_ _06239_ net528 vssd1 vssd1 vccd1 vccd1 _06240_ sky130_fd_sc_hd__mux2_1
X_11194_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[118\] _07104_
+ _07110_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[54\] _07152_
+ vssd1 vssd1 vccd1 vccd1 _07159_ sky130_fd_sc_hd__a221o_1
XFILLER_0_24_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11694__A team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[27\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13385__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17810_ clknet_leaf_91_wb_clk_i _03153_ _01506_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08582__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10145_ _04533_ net363 vssd1 vssd1 vccd1 vccd1 _06173_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17741_ clknet_leaf_91_wb_clk_i _03084_ _01437_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[51\]
+ sky130_fd_sc_hd__dfrtp_1
X_10076_ net895 _06104_ vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__nor2_1
X_14953_ net1215 vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__inv_2
XANTENNA__11981__X _07793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08334__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13904_ net1572 net981 _03788_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[23\]
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_89_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17672_ clknet_leaf_90_wb_clk_i _03015_ _01368_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[110\]
+ sky130_fd_sc_hd__dfrtp_1
X_14884_ net1230 vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16623_ clknet_leaf_141_wb_clk_i _02253_ _00319_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_950 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13835_ net1454 net579 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[13\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__12729__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_67_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08098__A1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16554_ clknet_leaf_195_wb_clk_i _02184_ _00250_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09611__B net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13766_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[17\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[16\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[19\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[18\]
+ vssd1 vssd1 vccd1 vccd1 _03739_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_139_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1008 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09295__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10978_ net961 _06481_ _06959_ vssd1 vssd1 vccd1 vccd1 _06960_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09834__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15505_ net1172 vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__inv_2
X_12717_ net302 net2832 net497 vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16485_ clknet_leaf_22_wb_clk_i _02115_ _00181_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13697_ team_05_WB.instance_to_wrap.wishbone.curr_state\[2\] _04169_ _07488_ team_05_WB.instance_to_wrap.wishbone.curr_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18224_ clknet_leaf_79_wb_clk_i net1455 _01919_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_15436_ net1164 vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12648_ net1003 _03686_ vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09047__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_84_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_155_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_154_Left_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09598__A1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18155_ clknet_leaf_0_wb_clk_i _03458_ _01851_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12464__S net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15367_ net1106 vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__inv_2
X_12579_ net500 net1857 net203 vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__mux2_1
XANTENNA__12317__X _03612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_152_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17106_ clknet_leaf_136_wb_clk_i _02736_ _00802_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_152_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14318_ net378 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[23\]
+ _04777_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__a22o_1
X_18086_ clknet_leaf_70_wb_clk_i _03409_ _01782_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[3\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold306 net79 vssd1 vssd1 vccd1 vccd1 net1720 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15298_ net1217 vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__inv_2
Xhold317 team_05_WB.instance_to_wrap.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 net1731
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[89\] vssd1 vssd1
+ vccd1 vccd1 net1742 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold339 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[3\] vssd1
+ vssd1 vccd1 vccd1 net1753 sky130_fd_sc_hd__dlygate4sd3_1
X_17037_ clknet_leaf_162_wb_clk_i _02667_ _00733_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_14249_ _04024_ _04034_ vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout808 net809 vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__buf_4
Xfanout819 net821 vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__clkbuf_8
X_08810_ net377 _04878_ vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__nand2b_2
XANTENNA__08573__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09790_ _05816_ _05820_ _05331_ vssd1 vssd1 vccd1 vccd1 _05821_ sky130_fd_sc_hd__a21bo_1
XANTENNA__12052__X _07864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10380__A2 _06390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1006 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net2420 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_163_Left_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1017 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2431 sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ _04806_ _04808_ _04810_ _04812_ vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__or4_2
X_17939_ clknet_leaf_35_wb_clk_i _03278_ _01635_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1028 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1039 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 net2453 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12212__B team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08325__A2 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08672_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[23\]
+ net816 net788 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_1032 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12639__S _03682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09286__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11632__A2 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1076_A net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_172_Left_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09224_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[10\]
+ net826 net778 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__a22o_1
XANTENNA__12374__S net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09155_ _04353_ _05209_ net954 vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12593__A0 _03612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1243_A net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08106_ net1032 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[8\]
+ net975 _04202_ vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09086_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[13\]
+ net591 _05137_ _05143_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[13\]
+ sky130_fd_sc_hd__o22a_4
XFILLER_0_71_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08037_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[13\] vssd1 vssd1
+ vccd1 vccd1 _04159_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1031_X net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold840 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold851 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net2265 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold862 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2276 sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net2287 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09210__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold884 team_05_WB.instance_to_wrap.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 net2298
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11699__A2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[24\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout870_A _04287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout491_X net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold895 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2309 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout968_A _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08564__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09988_ _06009_ _06016_ net526 vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__mux2_1
XANTENNA__10371__A2 _06387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_129_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_157_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08939_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[16\]
+ net837 net752 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[16\]
+ _05002_ vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_150_Right_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout756_X net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1540 team_05_WB.instance_to_wrap.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 net2954
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08316__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1551 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2965 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11950_ _07757_ _07760_ _07753_ _07756_ vssd1 vssd1 vccd1 vccd1 _07762_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_54_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10901_ _06895_ _06896_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[30\]
+ net565 vssd1 vssd1 vccd1 vccd1 _03436_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_93_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12549__S _03678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11881_ _07652_ _07659_ _07662_ vssd1 vssd1 vccd1 vccd1 _07693_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_28_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11453__S net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13620_ net1999 net328 net394 vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__mux2_1
X_10832_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[7\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06829_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_45_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09277__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09816__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13551_ net2074 net304 net402 vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10763_ _06759_ _06760_ net527 vssd1 vssd1 vccd1 vccd1 _06761_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_82_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12502_ net1639 _07821_ _03673_ vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16270_ net1115 vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__inv_2
XANTENNA__09029__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13482_ net289 net2964 net408 vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__mux2_1
X_10694_ net374 net361 _06120_ vssd1 vssd1 vccd1 vccd1 _06696_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15221_ net1061 vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__inv_2
X_12433_ net1657 _07816_ _03667_ vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15152_ net1185 vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__inv_2
X_12364_ _03607_ _03625_ _03630_ _03658_ vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__or4b_4
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14103_ _03968_ _03858_ _03967_ vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__or3b_1
XANTENNA_clkbuf_leaf_168_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11315_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[96\] _07123_
+ _07124_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[24\] _07273_
+ vssd1 vssd1 vccd1 vccd1 _07274_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15083_ net1068 vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__inv_2
XANTENNA__14325__B2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12295_ _03511_ _03589_ _03588_ _03586_ _03552_ vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__a2111o_1
X_14034_ _03874_ _03903_ vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__nand2b_1
X_11246_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[35\] _07097_
+ _07105_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[11\] vssd1 vssd1
+ vccd1 vccd1 _07208_ sky130_fd_sc_hd__a22o_1
XANTENNA__08555__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11177_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[127\] _07099_
+ _07124_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[31\] _07142_
+ vssd1 vssd1 vccd1 vccd1 _07143_ sky130_fd_sc_hd__a221o_1
XANTENNA__09606__B net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12639__A1 _07821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10128_ _06148_ _06155_ net530 vssd1 vssd1 vccd1 vccd1 _06156_ sky130_fd_sc_hd__mux2_1
X_15985_ net1140 vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08307__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17724_ clknet_leaf_86_wb_clk_i _03067_ _01420_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[34\]
+ sky130_fd_sc_hd__dfrtp_1
X_10059_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[7\] team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[6\]
+ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[5\] _06086_ vssd1 vssd1
+ vccd1 vccd1 _06088_ sky130_fd_sc_hd__and4_1
X_14936_ net1200 vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_29_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_106_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12459__S _03670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17655_ clknet_leaf_53_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[22\]
+ _01351_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_14867_ net1212 vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13818_ net1686 net971 net726 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[29\]
+ sky130_fd_sc_hd__and3_1
X_16606_ clknet_leaf_162_wb_clk_i _02236_ _00302_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_17586_ clknet_leaf_72_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[23\]
+ _01282_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09268__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14798_ net1184 vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16537_ clknet_leaf_9_wb_clk_i _02167_ _00233_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13749_ _05212_ _06464_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[17\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_154_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16468_ clknet_leaf_128_wb_clk_i _02098_ _00164_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14013__B1 _07451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18207_ clknet_leaf_38_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[28\]
+ _01902_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_15419_ net1123 vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16399_ clknet_leaf_135_wb_clk_i _02029_ _00095_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10707__S net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12575__A0 _03641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18138_ clknet_leaf_192_wb_clk_i _03441_ _01834_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold103 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[26\]
+ vssd1 vssd1 vccd1 vccd1 net1517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[25\]
+ vssd1 vssd1 vccd1 vccd1 net1528 sky130_fd_sc_hd__dlygate4sd3_1
X_18069_ clknet_leaf_95_wb_clk_i _03407_ _01765_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.lcd_rs
+ sky130_fd_sc_hd__dfrtp_1
Xhold125 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1539 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08794__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold136 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[21\]
+ vssd1 vssd1 vccd1 vccd1 net1550 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12922__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10008__A _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold147 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[17\]
+ vssd1 vssd1 vccd1 vccd1 net1561 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold158 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[23\]
+ vssd1 vssd1 vccd1 vccd1 net1572 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ net375 _05419_ vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__and2b_1
Xhold169 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[6\]
+ vssd1 vssd1 vccd1 vccd1 net1583 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout605 _04321_ vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__buf_4
XANTENNA__08546__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout616 _04318_ vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__buf_4
X_09842_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[20\]
+ net833 net806 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[20\]
+ _05872_ vssd1 vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__a221o_1
Xfanout627 net628 vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__buf_4
XFILLER_0_0_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout638 _04312_ vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__clkbuf_8
Xfanout649 net650 vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__clkbuf_8
XANTENNA__14141__C net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09773_ _05668_ _05803_ _05667_ vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__a21bo_2
X_08724_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[22\]
+ net593 _04787_ _04796_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[22\]
+ sky130_fd_sc_hd__o22a_2
X_08655_ _04724_ _04725_ _04726_ _04728_ vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__or4_1
XANTENNA__10510__C1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17522__Q team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[25\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout451_A _03714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11126__X _07092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout549_A _07448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08586_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[25\]
+ net839 net780 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout337_X net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout716_A _04286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09207_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[30\] _04246_
+ _04352_ _05258_ _05259_ vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__o311a_2
XFILLER_0_173_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09138_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[11\]
+ net682 net594 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09431__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08314__C net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08785__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09069_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[13\]
+ net810 net752 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__a22o_1
XANTENNA__12832__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11100_ _07065_ _07066_ vssd1 vssd1 vccd1 vccd1 _07067_ sky130_fd_sc_hd__nor2_1
X_12080_ _07888_ _07890_ _07884_ vssd1 vssd1 vccd1 vccd1 _07892_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold670 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2084 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout873_X net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold681 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[127\] vssd1 vssd1
+ vccd1 vccd1 net2095 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14332__B team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11448__S net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08537__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold692 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 net2106 sky130_fd_sc_hd__dlygate4sd3_1
X_11031_ net1046 _06669_ _07002_ net959 vssd1 vssd1 vccd1 vccd1 _07003_ sky130_fd_sc_hd__o211a_1
XANTENNA__13229__A team_05_WB.instance_to_wrap.total_design.core.instr_fetch vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08330__B net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13663__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15770_ net1297 vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09498__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12982_ net279 net2584 net464 vssd1 vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_86_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1370 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2784 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input12_A DAT_I[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1381 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2795 sky130_fd_sc_hd__dlygate4sd3_1
X_14721_ net1228 vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11933_ _07528_ _07744_ vssd1 vssd1 vccd1 vccd1 _07745_ sky130_fd_sc_hd__and2_1
XFILLER_0_169_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1392 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2806 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17440_ clknet_leaf_64_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[8\]
+ _01136_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_14652_ net1083 vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__inv_2
X_11864_ _07674_ _07675_ vssd1 vssd1 vccd1 vccd1 _07676_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13603_ net2423 net249 net394 vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__mux2_1
X_17371_ clknet_leaf_66_wb_clk_i net1445 _01067_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10815_ _06810_ _06811_ vssd1 vssd1 vccd1 vccd1 _06812_ sky130_fd_sc_hd__nor2_1
X_14583_ net1102 vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11795_ _07602_ _07603_ _07598_ _07599_ vssd1 vssd1 vccd1 vccd1 _07607_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_55_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16322_ net1139 vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_60_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13534_ net2275 net234 net402 vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10746_ net888 _06742_ _06744_ _05924_ vssd1 vssd1 vccd1 vccd1 _06745_ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16253_ net1133 vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_147_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_147_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13465_ net222 net2186 net410 vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10677_ net529 _06679_ net335 vssd1 vssd1 vccd1 vccd1 _06680_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15204_ net1229 vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__inv_2
X_12416_ _03610_ net1822 net214 vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__mux2_1
X_16184_ net1144 vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__inv_2
X_13396_ net2774 net193 net418 vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__mux2_1
XANTENNA__09422__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08776__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15135_ net1178 vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__inv_2
X_12347_ net545 _07507_ vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12742__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1086 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15066_ net1055 vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12278_ _07982_ _07983_ _07985_ _03570_ _03571_ vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__a2111o_1
X_14017_ _03864_ _03884_ _03886_ _03885_ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__a31o_1
XANTENNA__08528__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11229_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[4\] _07092_ _07101_
+ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[12\] _07191_ vssd1 vssd1
+ vccd1 vccd1 _07192_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10335__A2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08240__B net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13573__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15354__A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09489__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15968_ net1266 vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_125_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11296__B1 _07117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17707_ clknet_leaf_89_wb_clk_i _03050_ _01403_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[81\]
+ sky130_fd_sc_hd__dfrtp_1
X_14919_ net1104 vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__inv_2
X_15899_ net1301 vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08700__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08440_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[28\]
+ net646 net600 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[28\]
+ _04518_ vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__a221o_1
X_17638_ clknet_leaf_67_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[5\]
+ _01334_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_19_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08371_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[30\]
+ net838 net779 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12917__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17569_ clknet_leaf_113_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[6\]
+ _01265_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_173_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11599__B2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[25\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12548__A0 _03651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_3_0_wb_clk_i_X clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08767__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[21\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09964__A1 _04573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11220__B1 _07117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10574__A2 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09086__X team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08431__A _04510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17517__Q team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[20\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout402 net403 vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08519__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout413 _03727_ vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__clkbuf_4
Xfanout424 _03724_ vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__buf_8
XFILLER_0_10_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1206_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout435 _03722_ vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__clkbuf_4
Xfanout446 net447 vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__clkbuf_8
XANTENNA_input4_A DAT_I[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09825_ _05850_ _05852_ _05853_ _05855_ vssd1 vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__or4_2
XANTENNA__09192__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout457 _03712_ vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__clkbuf_4
Xfanout468 net471 vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__buf_6
XANTENNA_fanout666_A _04305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout479 _03705_ vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__buf_4
XANTENNA__13483__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09756_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[0\]
+ net648 net629 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__a22o_1
XANTENNA__11287__B1 _07125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08707_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[22\]
+ net834 net740 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[22\]
+ _04779_ vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09687_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[1\]
+ net707 net621 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout833_A net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout454_X net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08638_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[24\]
+ _04366_ net851 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[24\]
+ net856 vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_750 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08309__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout621_X net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08569_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[25\]
+ net701 net599 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[25\]
+ _04644_ vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__a221o_1
XANTENNA__12827__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout719_X net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10600_ _05820_ _05956_ _04279_ vssd1 vssd1 vccd1 vccd1 _06607_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_119_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11580_ net2477 net1006 _07392_ net358 vssd1 vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10531_ _06397_ _06503_ vssd1 vssd1 vccd1 vccd1 _06542_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10347__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12539__A0 _07836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13250_ net291 net2679 net437 vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__mux2_1
X_10462_ _06095_ _06476_ vssd1 vssd1 vccd1 vccd1 _06477_ sky130_fd_sc_hd__or2_1
XANTENNA__09404__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12201_ _07995_ _07998_ _07992_ vssd1 vssd1 vccd1 vccd1 _08013_ sky130_fd_sc_hd__a21o_1
XANTENNA__11211__B1 _07125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09955__A1 _05977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08758__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12562__S _03678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13181_ net293 net2380 net440 vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10393_ _06376_ _06410_ net520 vssd1 vssd1 vccd1 vccd1 _06411_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12132_ _07871_ _07891_ vssd1 vssd1 vccd1 vccd1 _07944_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_36_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12063_ _07524_ _07867_ _07536_ net543 vssd1 vssd1 vccd1 vccd1 _07875_ sky130_fd_sc_hd__a211o_1
X_16940_ clknet_leaf_1_wb_clk_i _02570_ _00636_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10317__A2 _06333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12711__A0 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11014_ _06619_ _06768_ _06898_ _06988_ net569 vssd1 vssd1 vccd1 vccd1 _06989_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_53_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16871_ clknet_leaf_203_wb_clk_i _02501_ _00567_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13393__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout980 team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[8\] vssd1 vssd1
+ vccd1 vccd1 net980 sky130_fd_sc_hd__buf_2
X_15822_ net1263 vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__inv_2
Xfanout991 _07481_ vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__buf_2
XANTENNA__08930__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15753_ net1295 vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_142_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12965_ net192 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[29\]
+ net465 vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_142_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09603__C net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14704_ net1093 vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11916_ _07702_ _07706_ _07727_ _07701_ vssd1 vssd1 vccd1 vccd1 _07728_ sky130_fd_sc_hd__o22a_1
X_15684_ net1156 vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ net196 net2114 net474 vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17423_ clknet_leaf_57_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[23\]
+ _01119_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_14635_ net1067 vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__inv_2
X_11847_ net549 _07657_ vssd1 vssd1 vccd1 vccd1 _07659_ sky130_fd_sc_hd__nand2_1
XANTENNA__12737__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17354_ clknet_leaf_38_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[18\]
+ _01050_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14566_ net1280 vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11778_ _07577_ _07578_ vssd1 vssd1 vccd1 vccd1 _07590_ sky130_fd_sc_hd__and2_1
XFILLER_0_144_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16305_ net1175 vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__inv_2
X_13517_ net2692 net294 net406 vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__mux2_1
X_17285_ clknet_leaf_176_wb_clk_i _02915_ _00981_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10729_ _05669_ _05803_ vssd1 vssd1 vccd1 vccd1 _06729_ sky130_fd_sc_hd__xor2_4
X_14497_ net1235 vssd1 vssd1 vccd1 vccd1 _00127_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16236_ net1136 vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload12 clknet_leaf_196_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload12/Y sky130_fd_sc_hd__clkinv_4
X_13448_ net2183 net290 net412 vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload23 clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload23/Y sky130_fd_sc_hd__inv_6
XFILLER_0_24_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload34 clknet_leaf_182_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload34/Y sky130_fd_sc_hd__clkinv_2
Xclkload45 clknet_leaf_194_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload45/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__08749__A2 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13568__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12472__S net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16167_ net1143 vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload56 clknet_leaf_179_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload56/Y sky130_fd_sc_hd__inv_6
XANTENNA__13795__C net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload67 clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload67/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_11_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13379_ net2193 net276 net422 vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__mux2_1
Xclkload78 clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload78/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_77_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload89 clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload89/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_149_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15118_ net1187 vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__inv_2
X_16098_ net1307 vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_149_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15049_ net1225 vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__inv_2
XFILLER_0_167_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09174__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08382__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09610_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[2\]
+ net877 net860 net857 vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__and4_1
XANTENNA__08921__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10720__S net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11269__B1 _07101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09541_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[3\]
+ net698 net676 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__a22o_1
XANTENNA__12995__X _03711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15812__A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09472_ _05512_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[4\]
+ sky130_fd_sc_hd__inv_2
X_08423_ _04494_ _04500_ _04501_ _04502_ vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__or4_2
XFILLER_0_65_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout247_A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08354_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[30\]
+ net645 net613 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10244__A1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[27\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08988__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload6 clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload6/Y sky130_fd_sc_hd__inv_8
XFILLER_0_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08285_ _04270_ _04347_ net945 net938 vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__o211a_4
XFILLER_0_6_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout414_A _03727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11992__A1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[25\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13986__B _07468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13478__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15259__A net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout202_X net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12382__S net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout783_A net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout210 net211 vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__buf_4
Xfanout1208 net1210 vssd1 vssd1 vccd1 vccd1 net1208 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1111_X net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1219 net1220 vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__buf_4
Xfanout221 _06248_ vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__clkbuf_2
Xfanout232 _06367_ vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09165__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout243 net244 vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout571_X net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout254 _06423_ vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__buf_2
XANTENNA_fanout950_A _04363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout265 net266 vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08373__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout669_X net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout276 net277 vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__clkbuf_2
X_09808_ _04970_ _05838_ _04967_ vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__a21oi_4
XANTENNA__08912__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout287 net289 vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__clkbuf_2
Xfanout298 _06621_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_4_15__f_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_15__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_09739_ net572 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[0\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[0\] vssd1 vssd1 vccd1
+ vccd1 _05770_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout836_X net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12750_ net298 net2052 net494 vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__mux2_1
X_11701_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[31\] team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[25\]
+ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[26\] team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[28\]
+ net993 vssd1 vssd1 vccd1 vccd1 _07513_ sky130_fd_sc_hd__o41a_1
XFILLER_0_96_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12557__S net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12681_ net2960 net342 vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__and2_1
XANTENNA__11461__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14420_ net1066 vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__inv_2
X_11632_ net107 net1012 _07354_ vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__a21o_1
XFILLER_0_139_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08979__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14351_ _04079_ _04069_ _04066_ _04065_ vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__o2bb2a_1
X_11563_ net1919 net1005 _07394_ net357 vssd1 vssd1 vccd1 vccd1 _03350_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13302_ net1944 net239 net430 vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__mux2_1
X_10514_ _06525_ vssd1 vssd1 vccd1 vccd1 _06526_ sky130_fd_sc_hd__inv_2
X_17070_ clknet_leaf_171_wb_clk_i _02700_ _00766_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14282_ _06572_ _06591_ _04055_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11494_ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[21\] net1003 vssd1
+ vssd1 vccd1 vccd1 _07405_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_98_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13388__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16021_ net1285 vssd1 vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__inv_2
XANTENNA__09928__A1 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15169__A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13233_ net219 net2793 net438 vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__mux2_1
X_10445_ _06457_ _06460_ vssd1 vssd1 vccd1 vccd1 _06461_ sky130_fd_sc_hd__or2_2
XFILLER_0_27_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_1068 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08600__A1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13164_ net219 net2513 net442 vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__mux2_1
X_10376_ _04778_ net367 _06043_ vssd1 vssd1 vccd1 vccd1 _06395_ sky130_fd_sc_hd__o21ai_1
X_12115_ _07923_ _07925_ _07921_ _07922_ vssd1 vssd1 vccd1 vccd1 _07927_ sky130_fd_sc_hd__a2bb2o_2
X_17972_ clknet_leaf_72_wb_clk_i _03311_ _01668_ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__dfrtp_1
X_13095_ net199 net2194 net450 vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__mux2_1
XANTENNA__10106__A _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09156__A2 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11499__B1 _07407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12046_ _07377_ _07468_ _07846_ vssd1 vssd1 vccd1 vccd1 _07858_ sky130_fd_sc_hd__or3_1
X_16923_ clknet_leaf_190_wb_clk_i _02553_ _00619_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_144_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08364__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16854_ clknet_leaf_141_wb_clk_i _02484_ _00550_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_161_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15805_ net1270 vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__inv_2
X_13997_ net978 team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[12\] vssd1
+ vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__nor2_1
X_16785_ clknet_leaf_172_wb_clk_i _02415_ _00481_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15736_ net1257 vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__inv_2
X_12948_ net283 net2657 net471 vssd1 vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10457__A2_N _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_162_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_162_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_34_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10474__A1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10474__B2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12467__S _03670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15667_ net1255 vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__inv_2
X_12879_ net274 net2431 net478 vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17406_ clknet_leaf_67_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[6\]
+ _01102_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14618_ net1055 vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__inv_2
X_18386_ net913 vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__clkbuf_1
X_15598_ net1258 vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17337_ clknet_leaf_39_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[1\]
+ _01033_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14549_ net1060 vssd1 vssd1 vccd1 vccd1 _00179_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08070_ net1024 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[26\]
+ net969 _04184_ vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11878__Y _07690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload101 clknet_leaf_153_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload101/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_70_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17268_ clknet_leaf_127_wb_clk_i _02898_ _00964_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload112 clknet_leaf_164_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload112/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_43_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload123 clknet_leaf_169_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload123/Y sky130_fd_sc_hd__bufinv_16
Xclkload134 clknet_leaf_144_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload134/Y sky130_fd_sc_hd__inv_6
XANTENNA__13298__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16219_ net1075 vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__inv_2
Xclkload145 clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload145/Y sky130_fd_sc_hd__clkinv_2
X_17199_ clknet_leaf_141_wb_clk_i _02829_ _00895_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload156 clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload156/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_113_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload167 clknet_leaf_85_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload167/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_168_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload178 clknet_leaf_110_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload178/X sky130_fd_sc_hd__clkbuf_8
Xclkload189 clknet_leaf_98_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload189/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__09395__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12930__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08972_ _05034_ vssd1 vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__inv_2
Xhold18 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[7\]
+ vssd1 vssd1 vccd1 vccd1 net1432 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[21\]
+ vssd1 vssd1 vccd1 vccd1 net1443 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08355__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10162__B1 _05924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10022__Y _06051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13100__A0 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout364_A _05770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09524_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[3\]
+ net810 net733 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09455_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[5\]
+ net740 _05490_ vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__a21o_1
XANTENNA__12377__S net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1273_A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout629_A _04314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08406_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[29\]
+ net665 _04485_ net720 vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__a211o_1
XFILLER_0_4_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09386_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[6\]
+ net615 net595 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_49_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08337_ net949 net938 _04418_ vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10768__A2 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout417_X net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08268_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[28\] team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[27\]
+ _04350_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__or3_1
XFILLER_0_50_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08199_ _04233_ net958 _04270_ _04152_ vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__a31o_1
XFILLER_0_85_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13001__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_35_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09386__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10230_ _06031_ _06040_ net530 vssd1 vssd1 vccd1 vccd1 _06255_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout786_X net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12390__A1 _03604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11193__A2 _07111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08594__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08322__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10161_ _05995_ _06187_ _05996_ net893 _05997_ vssd1 vssd1 vccd1 vccd1 _06188_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_7_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12840__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1005 net1006 vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__buf_2
XANTENNA__09138__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_58_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1016 _04347_ vssd1 vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__buf_1
Xfanout1027 net1030 vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__buf_2
XANTENNA__11964__B _07774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1038 net1039 vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_50_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10092_ net373 net366 vssd1 vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__and2_1
Xfanout1049 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write vssd1
+ vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__buf_4
XANTENNA__11456__S net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13920_ net1581 net981 _03796_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[31\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_96_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13851_ net1475 net578 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[29\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_88_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13671__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12802_ net241 net2486 net486 vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__mux2_1
X_13782_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[1\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[0\] team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[3\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[2\] vssd1
+ vssd1 vccd1 vccd1 _03755_ sky130_fd_sc_hd__or4_1
X_16570_ clknet_leaf_30_wb_clk_i _02200_ _00266_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10994_ net963 _06540_ _06972_ vssd1 vssd1 vccd1 vccd1 _06973_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10456__A1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15521_ net1154 vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12733_ net245 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[26\]
+ net495 vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__mux2_1
XANTENNA__09310__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15452_ net1149 vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__inv_2
X_18240_ clknet_leaf_66_wb_clk_i net1845 _01935_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_67_Left_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12664_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[25\]
+ net341 vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__and2_1
X_14403_ net1516 vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11979__X _07791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11615_ net112 net1011 net346 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[13\]
+ vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18171_ net1038 team_05_WB.instance_to_wrap.total_design.keypad0.next_rows\[3\] _01866_
+ vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__dfstp_1
XANTENNA_clkbuf_leaf_74_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15383_ net1103 vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__inv_2
X_12595_ _03645_ net2058 _03681_ vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_137_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13700__A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_756 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17122_ clknet_leaf_9_wb_clk_i _02752_ _00818_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_14334_ _04103_ _04104_ _04105_ _04106_ vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__or4_1
X_11546_ _07422_ _07425_ _07427_ net920 vssd1 vssd1 vccd1 vccd1 _07457_ sky130_fd_sc_hd__o31a_1
XFILLER_0_151_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18271__Q team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[25\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17053_ clknet_leaf_130_wb_clk_i _02683_ _00749_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_14265_ team_05_WB.instance_to_wrap.total_design.keypad0.counter\[3\] _04017_ vssd1
+ vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__or2_1
X_11477_ _07353_ _07387_ vssd1 vssd1 vccd1 vccd1 _07388_ sky130_fd_sc_hd__nor2_1
XANTENNA__12905__A0 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16004_ net1114 vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_74_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13216_ net298 net2362 net352 vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__mux2_1
X_10428_ _05972_ _06443_ net892 vssd1 vssd1 vccd1 vccd1 _06444_ sky130_fd_sc_hd__o21ai_1
X_14196_ _04000_ _04001_ net729 vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_164_Right_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11184__A2 _07097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12381__A1 _03614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08585__B1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_76_Left_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ net279 net2088 net444 vssd1 vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__mux2_1
X_10359_ _06161_ _06378_ net372 vssd1 vssd1 vccd1 vccd1 _06379_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12750__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10931__A2 _06918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09129__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ net272 net2864 net452 vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17955_ clknet_leaf_107_wb_clk_i _03294_ _01651_ vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09534__C1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12029_ _07363_ _07377_ vssd1 vssd1 vccd1 vccd1 _07841_ sky130_fd_sc_hd__or2_1
X_16906_ clknet_leaf_194_wb_clk_i _02536_ _00602_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_17886_ clknet_leaf_76_wb_clk_i _03229_ _01582_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_16837_ clknet_leaf_18_wb_clk_i _02467_ _00533_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13581__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10396__A2_N _06051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09837__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16768_ clknet_leaf_130_wb_clk_i _02398_ _00464_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10777__Y _06774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09301__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_85_Left_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15719_ net1142 vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16699_ clknet_leaf_189_wb_clk_i _02329_ _00395_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_18383__1368 vssd1 vssd1 vccd1 vccd1 _18383__1368/HI net1368 sky130_fd_sc_hd__conb_1
XFILLER_0_119_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09240_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[9\]
+ net706 net677 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__a22o_1
X_18391__1370 vssd1 vssd1 vccd1 vccd1 _18391__1370/HI net1370 sky130_fd_sc_hd__conb_1
XFILLER_0_29_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_926 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09171_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[11\]
+ net841 net790 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[11\]
+ _05224_ vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__a221o_1
X_18369_ net1354 vssd1 vssd1 vccd1 vccd1 la_data_out[17] sky130_fd_sc_hd__buf_2
XANTENNA__09065__A1 _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12925__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08122_ net1027 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[0\]
+ net969 _04210_ vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08053_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[5\] vssd1 vssd1
+ vccd1 vccd1 _04173_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09368__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_131_Right_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12372__A1 _07789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08576__B1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_119_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08955_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[15\]
+ net614 net606 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout481_A net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout579_A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08886_ _04950_ _04951_ vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09540__A2 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout746_A net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13491__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09507_ _05539_ _05541_ _05543_ _05545_ vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__or4_1
XFILLER_0_78_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout913_A net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08500__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10989__A2 _06521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09438_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[5\]
+ net674 net667 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[5\]
+ _05469_ vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__a221o_1
XFILLER_0_52_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09369_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[7\]
+ net851 net749 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[7\]
+ _05403_ vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout701_X net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12835__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11400_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[16\] _07330_
+ vssd1 vssd1 vccd1 vccd1 _07331_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12380_ net1619 _03620_ net217 vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11331_ net34 net35 net36 net37 vssd1 vssd1 vccd1 vccd1 _07289_ sky130_fd_sc_hd__or4b_2
XANTENNA__10610__A1 _06049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_895 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_158_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08333__B net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12348__D1 _07914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14050_ _03915_ _03917_ vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09359__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11262_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[43\] _07091_
+ _07099_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[123\] vssd1
+ vssd1 vccd1 vccd1 _07224_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_132_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11166__A2 _07100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13001_ net242 net2378 net463 vssd1 vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__mux2_1
XANTENNA__08567__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13666__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10213_ _06144_ _06154_ net518 vssd1 vssd1 vccd1 vccd1 _06239_ sky130_fd_sc_hd__mux2_1
X_11193_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[110\] _07111_
+ _07127_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[126\] _07157_
+ vssd1 vssd1 vccd1 vccd1 _07158_ sky130_fd_sc_hd__a221o_1
XANTENNA_input42_A wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10144_ net520 _06157_ _06171_ vssd1 vssd1 vccd1 vccd1 _06172_ sky130_fd_sc_hd__nand3_1
XFILLER_0_101_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17740_ clknet_leaf_93_wb_clk_i _03083_ _01436_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[50\]
+ sky130_fd_sc_hd__dfrtp_1
X_10075_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[31\] _06103_ vssd1
+ vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__xnor2_1
X_14952_ net1218 vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__inv_2
X_13903_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[23\]
+ net558 net577 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[23\]
+ net988 vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__a221o_1
X_17671_ clknet_leaf_76_wb_clk_i _03014_ _01367_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[109\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_89_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14883_ net1200 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__inv_2
X_16622_ clknet_leaf_169_wb_clk_i _02252_ _00318_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13834_ net1500 net579 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[12\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_98_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09819__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10597__Y _06605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18266__Q team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[20\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13765_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[21\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[20\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[23\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__or4_1
XFILLER_0_134_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16553_ clknet_leaf_14_wb_clk_i _02183_ _00249_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10977_ net1042 _06496_ _06958_ net956 vssd1 vssd1 vccd1 vccd1 _06959_ sky130_fd_sc_hd__o211a_1
XANTENNA__08098__A2 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09611__C net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15504_ net1166 vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__inv_2
X_12716_ net297 net2101 net498 vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__mux2_1
X_13696_ net1048 _06771_ _03689_ _03737_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.next_state\[1\]
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_clkbuf_leaf_197_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16484_ clknet_leaf_182_wb_clk_i _02114_ _00180_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18223_ clknet_leaf_79_wb_clk_i net1470 _01918_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13918__A2 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15435_ net1167 vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__inv_2
X_12647_ net1048 _06771_ vssd1 vssd1 vccd1 vccd1 _03686_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_156_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12745__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18154_ clknet_leaf_187_wb_clk_i _03457_ _01850_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_15366_ net1231 vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__inv_2
XANTENNA__09598__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12578_ _07859_ _07863_ _03659_ net919 vssd1 vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_124_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13787__D net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17105_ clknet_leaf_121_wb_clk_i _02735_ _00801_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11529_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[28\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[28\]
+ net1033 vssd1 vssd1 vccd1 vccd1 _07440_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_152_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14317_ net377 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[19\]
+ net376 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[18\] _04088_
+ vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__o221ai_2
XTAP_TAPCELL_ROW_152_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18085_ clknet_leaf_70_wb_clk_i _03408_ _01781_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_113_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15297_ net1225 vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold307 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[104\] vssd1 vssd1
+ vccd1 vccd1 net1721 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold318 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[93\] vssd1 vssd1
+ vccd1 vccd1 net1732 sky130_fd_sc_hd__dlygate4sd3_1
X_14248_ net2826 _04023_ vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__nor2_1
Xhold329 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[22\] vssd1 vssd1
+ vccd1 vccd1 net1743 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17036_ clknet_leaf_7_wb_clk_i _02666_ _00732_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13576__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12480__S _03673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14179_ team_05_WB.instance_to_wrap.CPU_DAT_O\[28\] net505 net909 vssd1 vssd1 vccd1
+ vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[28\] sky130_fd_sc_hd__and3_1
Xfanout809 _04391_ vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__buf_4
XFILLER_0_0_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08740_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[21\]
+ net608 net603 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[21\]
+ _04811_ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__a221o_1
Xhold1007 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 net2421 sky130_fd_sc_hd__dlygate4sd3_1
X_17938_ clknet_leaf_35_wb_clk_i _03277_ _01634_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1018 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 net2432 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2443 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09522__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08671_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[23\]
+ net847 net762 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[23\]
+ _04744_ vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__a221o_1
X_17869_ clknet_leaf_92_wb_clk_i _03212_ _01565_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08730__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18339__1328 vssd1 vssd1 vccd1 vccd1 _18339__1328/HI net1328 sky130_fd_sc_hd__conb_1
XFILLER_0_119_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09223_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[10\]
+ net840 net737 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[10\]
+ _05274_ vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__a221o_1
XFILLER_0_146_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout327_A _06753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1069_A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09154_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[30\] _04352_
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[20\] vssd1 vssd1
+ vccd1 vccd1 _05209_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_756 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09589__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08105_ net1032 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__and2b_1
XFILLER_0_115_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08797__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11131__Y _07097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14319__C1 _04091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09085_ _05139_ _05140_ _05141_ _05142_ vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__or4_1
XFILLER_0_130_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08036_ net1019 vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__inv_2
Xhold830 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2244 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold841 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2255 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13486__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08549__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout696_A net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold852 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 net2266 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12390__S _03660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold863 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold874 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net2288 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11699__A3 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[27\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold885 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net2310 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09761__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09987_ _06012_ _06015_ net512 vssd1 vssd1 vccd1 vccd1 _06016_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout484_X net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08938_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[16\]
+ net814 net741 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__a22o_1
Xhold1530 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net2944 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10659__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1541 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net2955 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1552 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 net2966 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout651_X net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08869_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[17\]
+ net620 _04318_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[17\]
+ _04935_ vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__a221o_1
XFILLER_0_99_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11320__A2 _07103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout749_X net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10900_ net960 _06108_ net565 vssd1 vssd1 vccd1 vccd1 _06896_ sky130_fd_sc_hd__a21o_1
XANTENNA__08721__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09712__B net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11880_ net549 _07690_ vssd1 vssd1 vccd1 vccd1 _07692_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_28_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10831_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[7\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06828_ sky130_fd_sc_hd__nand2_1
XANTENNA__18086__Q team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11608__B1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13550_ net2237 net296 net402 vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__mux2_1
X_10762_ _06113_ _06754_ net517 vssd1 vssd1 vccd1 vccd1 _06760_ sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12501_ net1663 _03666_ net210 vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13481_ net292 net2844 net408 vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__mux2_1
XANTENNA__12565__S net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10693_ _05552_ _06694_ net510 _05553_ vssd1 vssd1 vccd1 vccd1 _06695_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_54_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15220_ net1068 vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__inv_2
X_12432_ net1702 _07821_ _03667_ vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12033__B1 _07352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08344__A net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12584__A1 _07791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15151_ net1240 vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__inv_2
X_12363_ _03654_ _03655_ _03656_ _03657_ vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_130_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14102_ _03958_ _03961_ _03966_ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__o21a_1
X_11314_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[0\] _07092_ _07128_
+ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[64\] vssd1 vssd1 vccd1
+ vccd1 _07273_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_130_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15082_ net1121 vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__inv_2
X_12294_ _08008_ _03578_ _03582_ _03584_ vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__a31o_1
X_14033_ _03901_ _03902_ vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__or2_1
XANTENNA__13396__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11245_ net1877 net731 _07207_ vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18382__1367 vssd1 vssd1 vccd1 vccd1 _18382__1367/HI net1367 sky130_fd_sc_hd__conb_1
X_11176_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[95\] _07108_
+ _07123_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[103\] vssd1
+ vssd1 vccd1 vccd1 _07142_ sky130_fd_sc_hd__a22o_1
XANTENNA__09606__C net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08960__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10127_ _06151_ _06154_ net513 vssd1 vssd1 vccd1 vccd1 _06155_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15984_ net1141 vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__inv_2
XANTENNA__10114__A net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17723_ clknet_leaf_89_wb_clk_i _03066_ _01419_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09504__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10058_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[5\] _06086_ vssd1
+ vssd1 vccd1 vccd1 _06087_ sky130_fd_sc_hd__nand2_1
X_14935_ net1104 vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11311__A2 _07119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08712__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17654_ clknet_leaf_53_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[21\]
+ _01350_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_14866_ net1233 vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16605_ clknet_leaf_129_wb_clk_i _02235_ _00301_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13817_ net1587 net972 net724 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[28\]
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_158_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17585_ clknet_leaf_73_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[22\]
+ _01281_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_14797_ net1088 vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08238__B _04296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_69_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_85_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16536_ clknet_leaf_32_wb_clk_i _02166_ _00232_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_169_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13748_ net921 _06481_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[16\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11614__A3 _07472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16467_ clknet_leaf_166_wb_clk_i _02097_ _00163_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13798__C net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13679_ net2007 net293 net384 vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08491__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18206_ clknet_leaf_34_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[27\]
+ _01901_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_15418_ net1116 vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16398_ clknet_leaf_173_wb_clk_i _02028_ _00094_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_171_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08779__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18137_ clknet_leaf_11_wb_clk_i _03440_ _01833_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08243__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15349_ net1059 vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold104 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[23\]
+ vssd1 vssd1 vccd1 vccd1 net1518 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold115 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[6\]
+ vssd1 vssd1 vccd1 vccd1 net1529 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1000 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold126 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[30\]
+ vssd1 vssd1 vccd1 vccd1 net1540 sky130_fd_sc_hd__dlygate4sd3_1
X_18068_ clknet_leaf_99_wb_clk_i _03406_ _01764_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__dfrtp_1
Xhold137 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[4\]
+ vssd1 vssd1 vccd1 vccd1 net1551 sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1562 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold159 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[20\]
+ vssd1 vssd1 vccd1 vccd1 net1573 sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ _05350_ _05374_ vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17019_ clknet_leaf_191_wb_clk_i _02649_ _00715_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout606 _04320_ vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__clkbuf_8
X_09841_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[20\]
+ net752 net733 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05872_ sky130_fd_sc_hd__a22o_1
Xfanout617 net620 vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__clkbuf_8
Xfanout628 _04315_ vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__buf_4
XANTENNA__18398__A net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout639 _04312_ vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__clkbuf_4
XANTENNA__15815__A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09772_ _05734_ _05802_ _05733_ vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_28_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Left_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08723_ _04789_ _04791_ _04793_ _04795_ vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__or4_1
XANTENNA__10959__A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11302__A2 _07091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08654_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[23\]
+ net677 net670 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[23\]
+ _04727_ vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__a221o_1
XANTENNA__10311__X _06333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08585_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[25\]
+ net835 net816 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[25\]
+ _04658_ vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout444_A net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1186_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08467__C1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12385__S _07852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08482__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout611_A _04319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout709_A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09206_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[22\] net966
+ vssd1 vssd1 vccd1 vccd1 _05259_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_22_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08164__A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12566__A1 _07798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11369__A2 _06743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09137_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[11\]
+ net687 net656 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09068_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[13\]
+ net744 net737 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__a22o_1
XANTENNA__12318__A1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[18\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_898 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout699_X net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10633__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold660 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2074 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09707__B net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold671 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 net2085 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold682 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[55\] vssd1 vssd1
+ vccd1 vccd1 net2096 sky130_fd_sc_hd__dlygate4sd3_1
X_11030_ _06830_ _06831_ _06850_ _07001_ vssd1 vssd1 vccd1 vccd1 _07002_ sky130_fd_sc_hd__a31o_1
XANTENNA__09195__B1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold693 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2107 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09734__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout866_X net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08330__C net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12981_ net282 net2299 net465 vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_86_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11464__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1360 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2774 sky130_fd_sc_hd__dlygate4sd3_1
X_14720_ net1196 vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__inv_2
Xhold1371 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net2785 sky130_fd_sc_hd__dlygate4sd3_1
X_11932_ _07728_ _07743_ _07726_ vssd1 vssd1 vccd1 vccd1 _07744_ sky130_fd_sc_hd__o21ai_1
Xhold1382 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2796 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10501__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1393 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net2807 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08339__A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14651_ net1098 vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__inv_2
X_11863_ _07642_ _07643_ _07648_ _07635_ vssd1 vssd1 vccd1 vccd1 _07675_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10814_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[14\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06811_ sky130_fd_sc_hd__nor2_1
X_13602_ net2622 net227 net394 vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17370_ clknet_leaf_66_wb_clk_i net1422 _01066_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14582_ net1091 vssd1 vssd1 vccd1 vccd1 _00212_ sky130_fd_sc_hd__inv_2
X_11794_ _07605_ vssd1 vssd1 vccd1 vccd1 _07606_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16321_ net1132 vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_60_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13533_ net1997 net240 net403 vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__mux2_1
X_10745_ net888 _06743_ vssd1 vssd1 vccd1 vccd1 _06744_ sky130_fd_sc_hd__nand2_1
XANTENNA__08473__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16252_ net1140 vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__inv_2
XANTENNA__10280__A2 _06051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13464_ net220 net2245 net411 vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10676_ _06645_ _06678_ net516 vssd1 vssd1 vccd1 vccd1 _06679_ sky130_fd_sc_hd__mux2_1
X_12415_ _03655_ net1860 net215 vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__mux2_1
X_15203_ net1200 vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__inv_2
X_16183_ net1144 vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__inv_2
X_13395_ net1982 net198 net418 vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__mux2_1
XANTENNA__10109__A _05208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12346_ _03638_ _03639_ _03640_ vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__or3_4
X_15134_ net1054 vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_187_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_187_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_58_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15065_ net1051 vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_116_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_116_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12277_ _03570_ _03571_ vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14016_ net980 net979 vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__nand2b_1
XANTENNA__09186__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11228_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[116\] _07103_
+ _07130_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[100\] vssd1
+ vssd1 vccd1 vccd1 _07191_ sky130_fd_sc_hd__a22o_1
XANTENNA__09725__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18338__1327 vssd1 vssd1 vccd1 vccd1 _18338__1327/HI net1327 sky130_fd_sc_hd__conb_1
XFILLER_0_156_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08933__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08240__C net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11159_ _07039_ _07107_ vssd1 vssd1 vccd1 vccd1 _07125_ sky130_fd_sc_hd__nor2_4
XFILLER_0_156_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12611__X _03682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10740__B1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15967_ net1301 vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__inv_2
XFILLER_0_164_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17706_ clknet_leaf_95_wb_clk_i _03049_ _01402_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[80\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14918_ net1247 vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__inv_2
X_15898_ net1296 vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17637_ clknet_leaf_67_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[4\]
+ _01333_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_19_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14849_ net1236 vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11048__A1 _04170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08370_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[30\]
+ net834 net772 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[30\]
+ _04450_ vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__a221o_1
X_17568_ clknet_leaf_110_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[5\]
+ _01264_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_173_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16519_ clknet_leaf_202_wb_clk_i _02149_ _00215_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08464__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17499_ clknet_leaf_114_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[2\]
+ _01195_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_129_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12933__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14714__A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09177__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout403 _03730_ vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout414 _03727_ vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__buf_6
Xfanout425 _03724_ vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout394_A net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout436 _03721_ vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__buf_8
X_09824_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[20\]
+ net625 net606 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[20\]
+ _05854_ vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__a221o_1
Xfanout447 _03715_ vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__clkbuf_8
Xfanout458 _03712_ vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__buf_8
Xfanout469 net471 vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__buf_6
Xclkbuf_4_14__f_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_14__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09755_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[0\]
+ net880 net866 net863 vssd1 vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__and4_1
XANTENNA__11137__X _07103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08706_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[22\]
+ net828 net775 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__a22o_1
X_09686_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[1\]
+ net883 net871 net864 vssd1 vssd1 vccd1 vccd1 _05719_ sky130_fd_sc_hd__and4_1
XFILLER_0_68_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08637_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[24\]
+ net847 net807 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[24\]
+ _04701_ vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout826_A _04383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout447_X net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08568_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[25\]
+ net713 net678 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_Left_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09101__B1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18381__1366 vssd1 vssd1 vccd1 vccd1 _18381__1366/HI net1366 sky130_fd_sc_hd__conb_1
XFILLER_0_7_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08499_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[27\]
+ net775 net769 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout614_X net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08455__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13004__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10530_ net888 _06540_ _06539_ net554 vssd1 vssd1 vccd1 vccd1 _06541_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_36_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10461_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[17\] _06094_ vssd1
+ vssd1 vccd1 vccd1 _06476_ sky130_fd_sc_hd__nor2_1
XANTENNA__12843__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12200_ _07990_ _08011_ _07995_ vssd1 vssd1 vccd1 vccd1 _08012_ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09955__A2 _05978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13180_ net280 net2077 net441 vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__mux2_1
X_10392_ _06150_ _06152_ vssd1 vssd1 vccd1 vccd1 _06410_ sky130_fd_sc_hd__nand2_1
XANTENNA__08181__X _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11459__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12131_ _07881_ _07942_ vssd1 vssd1 vccd1 vccd1 _07943_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_36_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09168__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12062_ _07478_ _07870_ _07873_ vssd1 vssd1 vccd1 vccd1 _07874_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold490 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1904 sky130_fd_sc_hd__dlygate4sd3_1
X_11013_ _06854_ _06987_ vssd1 vssd1 vccd1 vccd1 _06988_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13674__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08915__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16870_ clknet_leaf_117_wb_clk_i _02500_ _00566_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10722__B1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout970 net973 vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__clkbuf_2
Xfanout981 net984 vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__clkbuf_4
X_15821_ net1256 vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__inv_2
Xfanout992 _07481_ vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_5_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15752_ net1257 vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__inv_2
X_12964_ net193 net2375 net466 vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09603__D net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09340__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1190 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2604 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_103_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14703_ net1283 vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__inv_2
X_11915_ _07707_ _07698_ vssd1 vssd1 vccd1 vccd1 _07727_ sky130_fd_sc_hd__and2b_1
X_15683_ net1156 vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ net197 net2633 net474 vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__mux2_1
XANTENNA__08694__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13262__X _03722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17422_ clknet_leaf_57_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[22\]
+ _01118_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13703__A net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14634_ net1110 vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__inv_2
X_11846_ _07657_ vssd1 vssd1 vccd1 vccd1 _07658_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17353_ clknet_leaf_37_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[17\]
+ _01049_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14565_ net1196 vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08446__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11777_ _07585_ _07588_ _07582_ vssd1 vssd1 vccd1 vccd1 _07589_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_166_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16304_ net1155 vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__inv_2
XANTENNA__11450__A1 _07346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13516_ net2520 net298 net405 vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__mux2_1
X_10728_ _05947_ _06727_ net888 vssd1 vssd1 vccd1 vccd1 _06728_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17284_ clknet_leaf_181_wb_clk_i _02914_ _00980_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14496_ net1195 vssd1 vssd1 vccd1 vccd1 _00126_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08235__C net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16235_ net1136 vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13447_ net2001 net278 net413 vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12753__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10659_ net515 _06127_ _06129_ _06662_ vssd1 vssd1 vccd1 vccd1 _06663_ sky130_fd_sc_hd__a31o_1
Xclkload13 clknet_leaf_197_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload13/Y sky130_fd_sc_hd__inv_8
XFILLER_0_23_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload24 clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload24/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_152_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload35 clknet_leaf_183_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload35/Y sky130_fd_sc_hd__bufinv_16
Xclkload46 clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload46/Y sky130_fd_sc_hd__bufinv_16
X_16166_ net1142 vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__inv_2
X_13378_ net2460 net272 net420 vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload57 clknet_leaf_180_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload57/X sky130_fd_sc_hd__clkbuf_8
Xclkload68 clknet_leaf_35_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload68/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_77_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload79 clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload79/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_77_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15117_ net1081 vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12329_ _03609_ _03619_ _03622_ _07774_ _03621_ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__a221o_1
X_16097_ net1307 vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_149_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15048_ net1223 vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08906__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13584__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_166_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10713__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16999_ clknet_leaf_201_wb_clk_i _02629_ _00695_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_84_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09540_ net570 net533 _05556_ vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__o21ai_4
XANTENNA__12212__A_N team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[14\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_13_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09471_ _04148_ _05510_ _05511_ vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__o21ba_1
X_08422_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[29\]
+ net840 net767 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[29\]
+ _04495_ vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08353_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[30\]
+ net618 net599 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__a22o_1
XANTENNA__08437__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10244__A2 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08284_ _04270_ net1017 net938 vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__o21a_4
XFILLER_0_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload7 clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload7/Y sky130_fd_sc_hd__inv_6
XFILLER_0_15_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1051_A net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14444__A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_25_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09538__A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10691__B net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17528__Q team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[31\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout200 _06107_ vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__clkbuf_2
Xfanout211 _03674_ vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13494__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout776_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1209 net1210 vssd1 vssd1 vccd1 vccd1 net1209 sky130_fd_sc_hd__buf_2
XANTENNA_fanout397_X net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout222 net225 vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__clkbuf_2
Xfanout233 _06367_ vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10911__S net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout244 net245 vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout255 _06442_ vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout266 _06462_ vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout277 _06537_ vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__clkbuf_2
X_09807_ _05014_ _05059_ _05836_ _05012_ vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__a31o_2
Xfanout288 net289 vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__buf_2
Xfanout299 _06621_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_105_Left_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09738_ net572 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[0\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[0\] vssd1 vssd1 vccd1
+ vccd1 _05769_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09322__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout731_X net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12838__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09669_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[1\]
+ net633 net598 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17640__D team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout829_X net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11700_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[26\] net995 vssd1
+ vssd1 vccd1 vccd1 _07512_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12680_ net2963 net341 vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__and2_1
XANTENNA__09720__B net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11631_ net1 _07344_ vssd1 vssd1 vccd1 vccd1 _07480_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_64_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_18337__1326 vssd1 vssd1 vccd1 vccd1 _18337__1326/HI net1326 sky130_fd_sc_hd__conb_1
XANTENNA__08428__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11562_ net93 net1004 net727 _07436_ vssd1 vssd1 vccd1 vccd1 _03351_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_145_Right_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14350_ _04082_ _04118_ _04120_ _04122_ vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__or4_1
XFILLER_0_52_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13669__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13301_ net2627 net242 net430 vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10513_ _06449_ _06524_ net528 vssd1 vssd1 vccd1 vccd1 _06525_ sky130_fd_sc_hd__mux2_1
X_14281_ _06609_ _06623_ _06641_ _04054_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__and4_1
X_11493_ _07346_ _07403_ vssd1 vssd1 vccd1 vccd1 _07404_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09389__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13232_ net191 net2716 net438 vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__mux2_1
X_16020_ net1285 vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input72_A wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10444_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[18\] net903 net966
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[18\] _06459_ vssd1
+ vssd1 vccd1 vccd1 _06460_ sky130_fd_sc_hd__a221o_1
XFILLER_0_150_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11196__B1 _07130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13163_ net189 net2910 net441 vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__mux2_1
X_10375_ net333 _06202_ _06207_ _06355_ _06393_ vssd1 vssd1 vccd1 vccd1 _06394_ sky130_fd_sc_hd__o221a_1
XFILLER_0_0_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08600__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[25\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12114_ _07923_ _07925_ vssd1 vssd1 vccd1 vccd1 _07926_ sky130_fd_sc_hd__nor2_1
X_17971_ clknet_leaf_73_wb_clk_i _03310_ _01667_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__dfrtp_1
X_13094_ _04257_ net563 _03695_ vssd1 vssd1 vccd1 vccd1 _03714_ sky130_fd_sc_hd__or3_4
XTAP_TAPCELL_ROW_72_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11499__A1 _07404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12045_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[31\] net1000 net543
+ vssd1 vssd1 vccd1 vccd1 _07857_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_72_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16922_ clknet_leaf_30_wb_clk_i _02552_ _00618_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_144_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_144_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16853_ clknet_leaf_22_wb_clk_i _02483_ _00549_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09614__C net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15804_ net1299 vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_161_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16784_ clknet_leaf_152_wb_clk_i _02414_ _00480_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10122__A _04818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13996_ _03862_ _03865_ vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09313__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15735_ net1301 vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12748__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12947_ net274 net2164 net470 vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__mux2_1
XANTENNA__08667__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15666_ net1257 vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__inv_2
X_12878_ net273 net2357 net476 vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__mux2_1
X_17405_ clknet_leaf_67_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[5\]
+ _01101_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14617_ net1052 vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__inv_2
X_18385_ net913 vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08419__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11829_ _07639_ _07640_ vssd1 vssd1 vccd1 vccd1 _07641_ sky130_fd_sc_hd__nand2_1
X_15597_ net1253 vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17336_ clknet_leaf_42_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[0\]
+ _01032_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14548_ net1074 vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09092__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13579__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12483__S _03673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17267_ clknet_leaf_168_wb_clk_i _02897_ _00963_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_131_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_131_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xclkload102 clknet_leaf_154_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload102/Y sky130_fd_sc_hd__clkinv_2
X_14479_ net1286 vssd1 vssd1 vccd1 vccd1 _00109_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload113 clknet_leaf_165_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload113/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_116_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload124 clknet_leaf_170_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload124/Y sky130_fd_sc_hd__bufinv_16
X_16218_ net1099 vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload135 clknet_leaf_145_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload135/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__08262__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[31\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17198_ clknet_leaf_175_wb_clk_i _02828_ _00894_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload146 clknet_leaf_130_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload146/Y sky130_fd_sc_hd__inv_6
Xclkload157 clknet_leaf_76_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload157/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__11187__B1 _07103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload168 clknet_leaf_86_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload168/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_168_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16149_ net1263 vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__inv_2
Xclkload179 clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload179/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_12_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08971_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[15\]
+ net715 _05024_ _05033_ vssd1 vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__o22a_4
XANTENNA_clkbuf_leaf_109_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold19 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[15\]
+ vssd1 vssd1 vccd1 vccd1 net1433 sky130_fd_sc_hd__dlygate4sd3_1
X_18380__1365 vssd1 vssd1 vccd1 vccd1 _18380__1365/HI net1365 sky130_fd_sc_hd__conb_1
XANTENNA__09552__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10032__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09523_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[3\]
+ net829 net822 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08658__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09454_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[5\]
+ net797 net750 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[5\]
+ _05495_ vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11134__Y _07100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08405_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[29\]
+ net694 net640 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__a22o_1
X_09385_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[6\]
+ net692 net645 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[6\]
+ _05428_ vssd1 vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__a221o_1
XFILLER_0_108_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08156__B net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08336_ _04236_ _04240_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[23\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[22\] _04230_ vssd1
+ vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__o2111a_2
XFILLER_0_117_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08724__X team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[22\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09083__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13489__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12393__S net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08267_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[26\] _04349_
+ vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_148_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_105_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08198_ _04232_ net962 _04271_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__o31a_1
XFILLER_0_21_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08172__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11178__B1 _07103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout893_A net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10160_ _05914_ _05927_ vssd1 vssd1 vccd1 vccd1 _06187_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout681_X net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08900__A team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[17\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1006 net1007 vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__clkbuf_2
XANTENNA__17635__D team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout779_X net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1017 _04347_ vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__clkbuf_4
X_10091_ net374 net361 _06118_ vssd1 vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__a21bo_1
XANTENNA__09715__B net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1028 net1030 vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_50_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1039 team_05_WB.instance_to_wrap.total_design.keypad0.key_clk vssd1 vssd1 vccd1
+ vccd1 net1039 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_50_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09543__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08897__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout946_X net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13890__A2 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13850_ net1482 net580 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[28\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_16_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12801_ net245 net2897 net486 vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__mux2_1
X_13781_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[5\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[4\] team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[7\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[6\] vssd1
+ vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__or4_1
X_10993_ _06551_ _06768_ _06898_ _06971_ net568 vssd1 vssd1 vccd1 vccd1 _06972_ sky130_fd_sc_hd__a221o_1
XANTENNA__08649__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11102__B1 _07031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15520_ net1154 vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__inv_2
X_12732_ net224 net2141 net494 vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_187_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15451_ net1149 vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09059__C1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12663_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[26\]
+ net342 vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__and2_1
X_14402_ net1529 vssd1 vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__clkbuf_1
X_18170_ net1038 team_05_WB.instance_to_wrap.total_design.keypad0.next_rows\[2\] _01865_
+ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__dfstp_1
XANTENNA__12602__A0 _03605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11614_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[14\] net997 _07472_
+ net1011 net2140 vssd1 vssd1 vccd1 vccd1 _03307_ sky130_fd_sc_hd__a32o_1
X_15382_ net1094 vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__inv_2
X_12594_ _03632_ net1775 net203 vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09074__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14355__Y _04128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17121_ clknet_leaf_149_wb_clk_i _02751_ _00817_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13399__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13700__B _06756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14333_ _05768_ _05801_ vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__nor2_1
X_11545_ net920 _07404_ _07405_ vssd1 vssd1 vccd1 vccd1 _07456_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08821__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17052_ clknet_leaf_157_wb_clk_i _02682_ _00748_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_162_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14264_ _04036_ _04043_ vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__nor2_1
X_11476_ net1001 _07386_ _07385_ vssd1 vssd1 vccd1 vccd1 _07387_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11169__B1 _07118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09609__C net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16003_ net1112 vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__inv_2
X_10427_ _04925_ _05933_ _05971_ vssd1 vssd1 vccd1 vccd1 _06443_ sky130_fd_sc_hd__and3_1
X_13215_ _06605_ net2952 net351 vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_74_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14195_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[3\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[4\]
+ _07027_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[5\] vssd1
+ vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10117__A _04989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13146_ net284 net2752 net447 vssd1 vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__mux2_1
X_10358_ _06283_ _06377_ net530 vssd1 vssd1 vccd1 vccd1 _06378_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13077_ net269 net2396 net452 vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__mux2_1
X_17954_ clknet_leaf_107_wb_clk_i _03293_ _01650_ vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_163_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10289_ _06297_ _06311_ _04275_ vssd1 vssd1 vccd1 vccd1 _06312_ sky130_fd_sc_hd__o21a_1
XANTENNA__10404__X _06422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12028_ _07794_ _07802_ _07808_ _07839_ vssd1 vssd1 vccd1 vccd1 _07840_ sky130_fd_sc_hd__or4b_4
XANTENNA__09534__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16905_ clknet_leaf_18_wb_clk_i _02535_ _00601_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_17885_ clknet_leaf_101_wb_clk_i _03228_ _01581_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08888__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16836_ clknet_leaf_184_wb_clk_i _02466_ _00532_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12478__S net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16767_ clknet_leaf_155_wb_clk_i _02397_ _00463_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13979_ _03848_ _03849_ vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__xor2_1
XFILLER_0_87_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15718_ net1142 vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16698_ clknet_leaf_11_wb_clk_i _02328_ _00394_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15649_ net1250 vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09170_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[11\]
+ net810 net760 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18368_ net1353 vssd1 vssd1 vccd1 vccd1 la_data_out[16] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_118_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08121_ net1027 net2305 vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__and2b_1
XFILLER_0_43_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17319_ clknet_leaf_200_wb_clk_i _02949_ _01015_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18299_ net1391 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
XANTENNA__13102__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08052_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[2\] vssd1 vssd1
+ vccd1 vccd1 _04172_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10027__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12941__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08954_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[15\]
+ net691 net602 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[15\]
+ _05016_ vssd1 vssd1 vccd1 vccd1 _05017_ sky130_fd_sc_hd__a221o_1
X_18336__1325 vssd1 vssd1 vccd1 vccd1 _18336__1325/HI net1325 sky130_fd_sc_hd__conb_1
XANTENNA__09525__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08885_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[17\]
+ net832 net771 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[17\]
+ _04948_ vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout474_A _03706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13625__X _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout641_A net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout262_X net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11145__X _07111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout739_A _04421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09506_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[4\]
+ net713 net696 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[4\]
+ _05544_ vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__a221o_1
XANTENNA__10438__A2 _06355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08167__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09437_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[5\]
+ net619 _05465_ net722 vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__a211o_1
XFILLER_0_94_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09368_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[7\]
+ net830 _05413_ net855 vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__a211o_1
XFILLER_0_47_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08454__X _04533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09056__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12060__A1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[11\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08319_ net942 net938 net935 vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09299_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[8\]
+ net662 _05347_ net722 vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__a211o_1
XANTENNA__08803__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13012__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11330_ net34 net37 net36 net35 vssd1 vssd1 vccd1 vccd1 _07288_ sky130_fd_sc_hd__or4b_1
XANTENNA__14337__B1 _05078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12348__C1 _07864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08333__C net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11261_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[75\] _07109_
+ _07111_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[107\] _07222_
+ vssd1 vssd1 vccd1 vccd1 _07223_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12851__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14632__A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13000_ net222 net2600 net462 vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__mux2_1
X_10212_ _06135_ _06147_ net518 vssd1 vssd1 vccd1 vccd1 _06238_ sky130_fd_sc_hd__mux2_1
X_11192_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[6\] _07092_ _07101_
+ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[14\] vssd1 vssd1 vccd1
+ vccd1 _07157_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10374__A1 _05887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10374__B2 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10143_ _04490_ net368 vssd1 vssd1 vccd1 vccd1 _06171_ sky130_fd_sc_hd__or2_1
XANTENNA_input35_A gpio_in[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10074_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[30\] team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[29\]
+ _06102_ vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__and3_1
X_14951_ net1242 vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11323__B1 _07116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13682__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13902_ net1569 net981 _03787_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[22\]
+ sky130_fd_sc_hd__o21a_1
X_17670_ clknet_leaf_78_wb_clk_i _03013_ _01366_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[108\]
+ sky130_fd_sc_hd__dfrtp_1
X_14882_ net1226 vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__inv_2
X_16621_ clknet_leaf_160_wb_clk_i _02251_ _00317_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13833_ net1483 net581 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[11\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_69_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16552_ clknet_leaf_204_wb_clk_i _02182_ _00248_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13764_ _04171_ net1884 net1031 vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11626__B2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10976_ _04170_ _06866_ _06957_ vssd1 vssd1 vccd1 vccd1 _06958_ sky130_fd_sc_hd__or3_1
XANTENNA__09295__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09611__D net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15503_ net1166 vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_139_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12715_ net300 net2230 net497 vssd1 vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16483_ clknet_leaf_198_wb_clk_i _02113_ _00179_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13695_ _06770_ net1048 vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__and2b_1
XFILLER_0_31_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18222_ clknet_leaf_79_wb_clk_i net1565 _01917_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15434_ net1158 vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__inv_2
X_12646_ team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.state\[1\] team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.state\[0\]
+ net1048 vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__or3b_1
XFILLER_0_26_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09047__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18153_ clknet_leaf_17_wb_clk_i _03456_ _01849_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08255__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15365_ net1193 vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__inv_2
X_12577_ _07850_ _03669_ _07840_ vssd1 vssd1 vccd1 vccd1 _03680_ sky130_fd_sc_hd__and3b_4
X_17104_ clknet_leaf_167_wb_clk_i _02734_ _00800_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14316_ net377 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__nor2_1
X_11528_ _07431_ _07434_ _07436_ _07438_ vssd1 vssd1 vccd1 vccd1 _07439_ sky130_fd_sc_hd__or4_1
X_18084_ clknet_leaf_83_wb_clk_i _00011_ _01780_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_152_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15296_ net1102 vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__inv_2
XANTENNA__12046__B _07468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold308 net86 vssd1 vssd1 vccd1 vccd1 net1722 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold319 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[85\] vssd1 vssd1
+ vccd1 vccd1 net1733 sky130_fd_sc_hd__dlygate4sd3_1
X_17035_ clknet_leaf_188_wb_clk_i _02665_ _00731_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_14247_ net1918 _04024_ vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__xor2_1
XANTENNA__12761__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11459_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[6\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[6\]
+ net1034 vssd1 vssd1 vccd1 vccd1 _07370_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14178_ net1624 net502 net908 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[27\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__11377__S net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13129_ net194 net2643 net445 vssd1 vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1008 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 net2422 sky130_fd_sc_hd__dlygate4sd3_1
X_17937_ clknet_leaf_34_wb_clk_i _03276_ _01633_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11314__B1 _07128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1019 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2433 sky130_fd_sc_hd__dlygate4sd3_1
X_08670_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[23\]
+ net799 net742 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12212__D team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17868_ clknet_leaf_84_wb_clk_i _03211_ _01564_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16819_ clknet_leaf_170_wb_clk_i _02449_ _00515_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17799_ clknet_leaf_89_wb_clk_i _03142_ _01495_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[109\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09286__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12936__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09222_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[10\]
+ net832 net736 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12508__Y _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09153_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[11\]
+ net715 _05202_ _05207_ vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__o22a_4
XANTENNA__12042__A1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[27\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08246__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08104_ net1030 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[9\]
+ net974 _04201_ vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__a22o_1
XANTENNA__14319__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09084_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[13\]
+ net822 net782 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[13\]
+ _05129_ vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__a221o_1
XFILLER_0_114_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08153__C team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08035_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[13\] vssd1
+ vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__inv_2
XANTENNA__15548__A net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold820 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 net2234 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_82_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold831 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net2245 sky130_fd_sc_hd__dlygate4sd3_1
Xhold842 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2256 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1229_A net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold853 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net2267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold864 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 net2278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold875 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2289 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09210__A2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout591_A _04368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold886 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 net2300 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout689_A net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold897 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 net2311 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10191__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09986_ _06013_ _06014_ vssd1 vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1017_X net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08937_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[16\]
+ net845 net806 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[16\]
+ _05000_ vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout477_X net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout856_A _04367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1520 net109 vssd1 vssd1 vccd1 vccd1 net2934 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1531 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 net2945 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1542 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 net2956 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1553 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 net2967 sky130_fd_sc_hd__dlygate4sd3_1
X_08868_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[17\]
+ net682 _04314_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09712__C net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08799_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[19\]
+ net830 net790 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[19\]
+ _04868_ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout644_X net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13007__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10830_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[8\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[8\]
+ vssd1 vssd1 vccd1 vccd1 _06827_ sky130_fd_sc_hd__nand2_1
XANTENNA__11608__A1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[17\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11608__B2 net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09277__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08485__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout811_X net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12846__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10761_ net512 _06723_ vssd1 vssd1 vccd1 vccd1 _06759_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout909_X net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12500_ net1633 _03665_ _03674_ vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10692_ net1020 _05551_ net552 vssd1 vssd1 vccd1 vccd1 _06694_ sky130_fd_sc_hd__a21oi_1
X_13480_ net280 net2825 net409 vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09029__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12431_ _03666_ net1799 net214 vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10366__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08344__B team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[31\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15150_ net1191 vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__inv_2
X_12362_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[25\] net1000 _03596_
+ _03626_ net543 vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__a2111o_4
X_14101_ _03958_ _03961_ _03966_ vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_130_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13677__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11313_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[88\] _07096_
+ _07111_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[104\] vssd1
+ vssd1 vccd1 vccd1 _07272_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12581__S net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12293_ _03578_ _03579_ _03587_ _03511_ vssd1 vssd1 vccd1 vccd1 _03588_ sky130_fd_sc_hd__o211a_1
X_15081_ net1225 vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11244_ _07194_ _07200_ _07206_ vssd1 vssd1 vccd1 vccd1 _07207_ sky130_fd_sc_hd__or3_1
X_14032_ _03866_ _03871_ _03900_ vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__and3_1
XANTENNA__09201__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11175_ _07077_ _07136_ _07138_ _07140_ vssd1 vssd1 vccd1 vccd1 _07141_ sky130_fd_sc_hd__or4_1
XANTENNA__09606__D net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10126_ _06152_ _06153_ vssd1 vssd1 vccd1 vccd1 _06154_ sky130_fd_sc_hd__nand2_1
X_15983_ net1141 vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17722_ clknet_leaf_95_wb_clk_i _03065_ _01418_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13706__A net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10057_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[4\] team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[3\]
+ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[2\] vssd1 vssd1 vccd1
+ vccd1 _06086_ sky130_fd_sc_hd__and3_1
X_14934_ net1085 vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_69_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18277__Q team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[31\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17653_ clknet_leaf_39_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[20\]
+ _01349_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_14865_ net1192 vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload0_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16604_ clknet_leaf_157_wb_clk_i _02234_ _00300_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13816_ net1492 net970 net723 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[27\]
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_158_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17584_ clknet_leaf_72_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[21\]
+ _01280_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09268__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14796_ net1109 vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_158_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16535_ clknet_leaf_146_wb_clk_i _02165_ _00231_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08238__C net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13747_ net921 _06500_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[15\]
+ sky130_fd_sc_hd__nor2_1
X_10959_ net956 _06424_ vssd1 vssd1 vccd1 vccd1 _06944_ sky130_fd_sc_hd__nor2_1
XANTENNA__12756__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16466_ clknet_leaf_120_wb_clk_i _02096_ _00162_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13678_ net2048 net281 net384 vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__mux2_1
XANTENNA__14013__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12328__Y _03623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18205_ clknet_leaf_35_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[26\]
+ _01900_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18335__1324 vssd1 vssd1 vccd1 vccd1 _18335__1324/HI net1324 sky130_fd_sc_hd__conb_1
XFILLER_0_128_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15417_ net1123 vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_2__f_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12629_ _03645_ net1903 net201 vssd1 vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__mux2_1
X_16397_ clknet_leaf_161_wb_clk_i _02027_ _00093_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_171_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_171_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_38_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_18136_ clknet_leaf_12_wb_clk_i _03439_ _01832_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15348_ net1068 vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09440__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13587__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12491__S net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18067_ clknet_leaf_103_wb_clk_i _03405_ _01763_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold105 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[16\]
+ vssd1 vssd1 vccd1 vccd1 net1519 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold116 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[26\]
+ vssd1 vssd1 vccd1 vccd1 net1530 sky130_fd_sc_hd__dlygate4sd3_1
X_15279_ net1286 vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__inv_2
Xhold127 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[4\]
+ vssd1 vssd1 vccd1 vccd1 net1541 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold138 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[16\]
+ vssd1 vssd1 vccd1 vccd1 net1552 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[0\]
+ vssd1 vssd1 vccd1 vccd1 net1563 sky130_fd_sc_hd__dlygate4sd3_1
X_17018_ clknet_leaf_11_wb_clk_i _02648_ _00714_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_1000 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08270__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[30\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09840_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[20\]
+ net822 net745 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[20\]
+ _05870_ vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__a221o_1
Xfanout607 _04320_ vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout618 net620 vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08400__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout629 _04314_ vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_13__f_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_13__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_09771_ net362 _05801_ vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__and2_2
XFILLER_0_119_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08722_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[22\]
+ net849 net809 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[22\]
+ _04794_ vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__a221o_1
XANTENNA__10959__B _06424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08653_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[23\]
+ net626 net608 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__a22o_1
XANTENNA__10510__A1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08584_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[25\]
+ net796 net739 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__a22o_1
XFILLER_0_166_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1081_A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout437_A _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11142__Y _07108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09205_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[30\] _05257_
+ vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_40_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12015__A1 _07478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13212__A0 _06554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout604_A net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09136_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[11\]
+ net644 net636 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09431__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13497__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09067_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[25\] net966
+ net955 _05125_ _04345_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[13\]
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold650 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net2064 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout973_A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold661 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net2075 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout594_X net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09707__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold672 net77 vssd1 vssd1 vccd1 vccd1 net2086 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold683 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 net2097 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold694 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2108 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09969_ _04491_ _04511_ _05996_ _05997_ vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout761_X net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout859_X net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09723__B net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12980_ net274 net2637 net467 vssd1 vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__mux2_1
XANTENNA__09498__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1350 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2764 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_86_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1361 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net2775 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_86_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11931_ _07730_ _07739_ _07742_ vssd1 vssd1 vccd1 vccd1 _07743_ sky130_fd_sc_hd__and3_1
Xhold1372 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2786 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10221__Y _06247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1383 team_05_WB.instance_to_wrap.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 net2797
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1394 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net2808 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08339__B net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14650_ net1055 vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11862_ _07644_ _07647_ vssd1 vssd1 vccd1 vccd1 _07674_ sky130_fd_sc_hd__or2_1
XFILLER_0_169_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13601_ net2030 net230 net394 vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__mux2_1
X_10813_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[14\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06810_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_0_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14581_ net1060 vssd1 vssd1 vccd1 vccd1 _00211_ sky130_fd_sc_hd__inv_2
XANTENNA__08458__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11793_ _07602_ _07603_ vssd1 vssd1 vccd1 vccd1 _07605_ sky130_fd_sc_hd__nor2_1
XANTENNA__11480__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16320_ net1131 vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__inv_2
XANTENNA__10265__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13532_ net1987 net243 net403 vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10744_ _05735_ _05802_ vssd1 vssd1 vccd1 vccd1 _06743_ sky130_fd_sc_hd__xor2_4
XFILLER_0_171_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16251_ net1132 vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_11_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13203__A0 _06384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13463_ net190 net2126 net408 vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__mux2_1
X_10675_ _06011_ _06013_ vssd1 vssd1 vccd1 vccd1 _06678_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15202_ net1226 vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__inv_2
X_12414_ _03646_ net1838 net215 vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16182_ net1144 vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__inv_2
X_13394_ net557 _03697_ _03701_ vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__and3_4
XANTENNA__09422__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15133_ net1087 vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__inv_2
X_12345_ _03531_ _03536_ vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08630__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13200__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15064_ net1207 vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12276_ _07978_ _03564_ _03566_ vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__and3_1
XANTENNA__11517__B1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09617__C net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14015_ net979 _03864_ vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__nor2_1
X_11227_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[92\] _07096_
+ _07127_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[124\] vssd1
+ vssd1 vccd1 vccd1 _07190_ sky130_fd_sc_hd__a22o_1
XANTENNA__10125__A net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11158_ _07087_ _07122_ vssd1 vssd1 vccd1 vccd1 _07124_ sky130_fd_sc_hd__nor2_4
Xclkbuf_leaf_156_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_156_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_147_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10740__A1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10109_ _05208_ net365 vssd1 vssd1 vccd1 vccd1 _06137_ sky130_fd_sc_hd__or2_1
X_11089_ _07032_ _07044_ _07055_ vssd1 vssd1 vccd1 vccd1 _07056_ sky130_fd_sc_hd__nand3_1
X_15966_ net1278 vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__inv_2
XANTENNA__09633__B net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09489__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17705_ clknet_leaf_99_wb_clk_i _03048_ _01401_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[79\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14917_ net1185 vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__inv_2
XANTENNA__11296__A2 _07115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12493__A1 _07812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15897_ net1275 vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_159_Right_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09920__Y _05949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17636_ clknet_leaf_70_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[3\]
+ _01332_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_14848_ net1195 vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12486__S net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08449__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17567_ clknet_leaf_113_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[4\]
+ _01263_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_14779_ net1099 vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08536__Y _04613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09110__A1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[24\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16518_ clknet_leaf_117_wb_clk_i _02148_ _00214_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17498_ clknet_leaf_114_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[1\]
+ _01194_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_105_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09661__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16449_ clknet_leaf_150_wb_clk_i _02079_ _00145_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18119_ clknet_leaf_45_wb_clk_i _00033_ _01815_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15098__A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11220__A2 _07115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13110__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10306__Y _06328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout404 net407 vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__buf_6
XFILLER_0_100_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14730__A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout415 _03727_ vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__buf_4
Xfanout426 _03724_ vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__buf_6
X_09823_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[20\]
+ net707 net676 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__a22o_1
Xfanout437 _03721_ vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__clkbuf_4
Xfanout448 _03714_ vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__buf_6
Xfanout459 _03712_ vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__buf_4
X_09754_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[0\]
+ net881 _04283_ net863 vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__and4_1
XANTENNA__10689__B _05807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08705_ _04777_ vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__inv_2
XANTENNA__11287__A2 _07104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12484__A1 _03646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08688__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09685_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[1\]
+ net876 net864 net860 vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout554_A net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_169_Left_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08636_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[24\]
+ net803 net754 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[24\]
+ _04698_ vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__a221o_1
XFILLER_0_68_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08567_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[25\]
+ net688 net615 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[25\]
+ _04642_ vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout721_A _04285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout342_X net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_54_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout819_A net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1000 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08498_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[27\]
+ net847 net734 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[27\]
+ _04575_ vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08175__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[11\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08860__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout607_X net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10460_ _06466_ _06474_ net536 vssd1 vssd1 vccd1 vccd1 _06475_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09404__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17638__D team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[5\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09119_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[12\]
+ net759 net737 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[12\]
+ _05174_ vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__a221o_1
XFILLER_0_161_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11211__A2 _07111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10391_ net892 _06408_ _06407_ _05924_ vssd1 vssd1 vccd1 vccd1 _06409_ sky130_fd_sc_hd__o211a_1
XANTENNA__08612__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_1__f_wb_clk_i_X clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13020__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12130_ _07871_ _07891_ vssd1 vssd1 vccd1 vccd1 _07942_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12061_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[11\] team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[12\]
+ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[13\] net998 net543 vssd1
+ vssd1 vccd1 vccd1 _07873_ sky130_fd_sc_hd__a41o_1
Xhold480 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[89\] vssd1 vssd1
+ vccd1 vccd1 net1894 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold491 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[24\] vssd1 vssd1
+ vccd1 vccd1 net1905 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11012_ _06825_ _06826_ vssd1 vssd1 vccd1 vccd1 _06987_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_53_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11475__S net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout960 net961 vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__buf_2
X_15820_ net1293 vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__inv_2
X_18334__1323 vssd1 vssd1 vccd1 vccd1 _18334__1323/HI net1323 sky130_fd_sc_hd__conb_1
Xfanout971 net973 vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__buf_2
Xfanout982 net984 vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__buf_2
Xfanout993 net994 vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_93_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15751_ net1292 vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__inv_2
XANTENNA__11278__A2 _07120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12963_ net197 net2870 net466 vssd1 vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__mux2_1
XANTENNA__08679__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1180 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net2594 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13690__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14702_ net1189 vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__inv_2
Xhold1191 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net2605 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11914_ _07725_ _07702_ _07703_ vssd1 vssd1 vccd1 vccd1 _07726_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15682_ net1148 vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__inv_2
X_12894_ _04253_ net562 _03702_ vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__or3_4
XTAP_TAPCELL_ROW_16_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ clknet_leaf_58_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[21\]
+ _01117_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14633_ net1221 vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__inv_2
X_18349__1334 vssd1 vssd1 vccd1 vccd1 _18349__1334/HI net1334 sky130_fd_sc_hd__conb_1
XANTENNA__13703__B _06706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11845_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[4\] net997 vssd1
+ vssd1 vccd1 vccd1 _07657_ sky130_fd_sc_hd__nand2_2
XANTENNA__11063__X _07030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17352_ clknet_leaf_37_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[16\]
+ _01048_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_14564_ net1232 vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11776_ _07587_ _07586_ _07584_ vssd1 vssd1 vccd1 vccd1 _07588_ sky130_fd_sc_hd__or3b_2
XFILLER_0_32_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16303_ net1155 vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13515_ net2432 net286 net407 vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__mux2_1
X_17283_ clknet_leaf_199_wb_clk_i _02913_ _00979_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10727_ _05669_ _05946_ vssd1 vssd1 vccd1 vccd1 _06727_ sky130_fd_sc_hd__or2_1
X_14495_ net1178 vssd1 vssd1 vccd1 vccd1 _00125_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08851__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16234_ net1136 vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09909__A _05256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13446_ net2301 net283 net413 vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09779__A_N _05442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10658_ net515 _06661_ vssd1 vssd1 vccd1 vccd1 _06662_ sky130_fd_sc_hd__nor2_1
Xclkload14 clknet_leaf_198_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload14/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_141_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_200_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkload25 clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload25/Y sky130_fd_sc_hd__inv_6
XFILLER_0_141_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16165_ net1142 vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__inv_2
Xclkload36 clknet_leaf_185_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload36/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_106_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13377_ net2941 net268 net420 vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__mux2_1
Xclkload47 clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload47/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload58 clknet_leaf_181_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload58/Y sky130_fd_sc_hd__clkinv_2
X_10589_ _06064_ _06596_ net332 _06450_ vssd1 vssd1 vccd1 vccd1 _06597_ sky130_fd_sc_hd__o2bb2a_1
Xclkload69 clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload69/Y sky130_fd_sc_hd__inv_4
XTAP_TAPCELL_ROW_77_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15116_ net1109 vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__inv_2
X_12328_ _07774_ _03622_ vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__nand2_4
XFILLER_0_11_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16096_ net1307 vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_149_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15047_ net1106 vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__inv_2
X_12259_ _07959_ _03553_ vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_166_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08382__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16998_ clknet_leaf_118_wb_clk_i _02628_ _00694_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11269__A2 _07092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12466__A1 _03666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15949_ net1270 vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__inv_2
X_09470_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[16\] net965
+ _04268_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[11\] _05354_
+ vssd1 vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08421_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[29\]
+ net833 _04497_ vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__a21o_1
X_17619_ clknet_leaf_58_wb_clk_i _02990_ _01315_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13105__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_53_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08352_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[30\]
+ net697 net673 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[30\]
+ _04430_ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09095__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08283_ _04150_ _04151_ _04237_ _04241_ _04231_ vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__a221o_1
XANTENNA__08842__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12944__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload8 clknet_leaf_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload8/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_138_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_74_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout302_A _06655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1044_A net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10952__A1 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1211_A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout201 _03683_ vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__buf_4
XFILLER_0_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout212 net213 vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__buf_4
XFILLER_0_10_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout223 net225 vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout234 net237 vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__clkbuf_2
Xfanout245 _06294_ vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__buf_2
Xfanout256 _06442_ vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_31_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout769_A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout267 net268 vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_31_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08373__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09806_ _05059_ _05836_ vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__nand2_2
XFILLER_0_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout278 net281 vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__buf_2
Xfanout289 _06606_ vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_2_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12457__A1 _03645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09737_ _05768_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[0\]
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_2_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout936_A net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09668_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[1\]
+ net878 net874 net869 vssd1 vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__and4_1
XFILLER_0_55_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_177_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08619_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[24\]
+ net645 net603 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[24\]
+ _04679_ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout724_X net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09720__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09599_ net571 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[2\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[2\] vssd1 vssd1 vccd1
+ vccd1 _05634_ sky130_fd_sc_hd__a21o_2
XANTENNA__13015__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11630_ net108 net1008 net345 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__a22o_1
XANTENNA__09625__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11561_ net1850 net1004 net727 _07409_ vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__a22o_1
XANTENNA__12854__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11611__X _07476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13300_ net2350 net223 net429 vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10512_ net513 _06143_ _06145_ _06523_ vssd1 vssd1 vccd1 vccd1 _06524_ sky130_fd_sc_hd__a31o_1
X_14280_ _06658_ _06672_ _06691_ _04053_ vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__and4_1
X_11492_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[21\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[21\]
+ net1031 vssd1 vssd1 vccd1 vccd1 _07403_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_98_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13231_ net193 net2480 net439 vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__mux2_1
X_10443_ net896 _06458_ vssd1 vssd1 vccd1 vccd1 _06459_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input65_A wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13162_ net195 net2787 net443 vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__mux2_1
X_10374_ _05887_ net510 _06210_ net337 _06392_ vssd1 vssd1 vccd1 vccd1 _06393_ sky130_fd_sc_hd__o221a_1
XFILLER_0_27_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13685__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12113_ _07914_ _07919_ vssd1 vssd1 vccd1 vccd1 _07925_ sky130_fd_sc_hd__xor2_1
X_17970_ clknet_leaf_105_wb_clk_i _03309_ _01666_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__dfrtp_1
X_13093_ net307 net1956 net453 vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12044_ _07508_ _07853_ _07854_ _07855_ vssd1 vssd1 vccd1 vccd1 _07856_ sky130_fd_sc_hd__or4_2
X_16921_ clknet_leaf_12_wb_clk_i _02551_ _00617_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09010__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08364__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09561__B2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16852_ clknet_leaf_115_wb_clk_i _02482_ _00548_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09614__D net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout790 net793 vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__clkbuf_8
X_15803_ net1302 vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_161_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12448__A1 _07793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16783_ clknet_leaf_134_wb_clk_i _02413_ _00479_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13995_ _03862_ _03863_ _03864_ vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__nand3_1
XFILLER_0_172_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13714__A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15734_ net1295 vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12946_ net271 net2764 net468 vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15665_ net1257 vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__inv_2
X_12877_ net267 net2878 net476 vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17404_ clknet_leaf_67_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[4\]
+ _01100_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_14616_ net1207 vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__inv_2
X_18384_ net913 vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09077__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11828_ _07576_ _07596_ _07559_ vssd1 vssd1 vccd1 vccd1 _07640_ sky130_fd_sc_hd__or3b_2
X_15596_ net1167 vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12049__B _07468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17335_ clknet_leaf_143_wb_clk_i _02965_ _01031_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14547_ net1216 vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__inv_2
XANTENNA__12620__A1 _07793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11759_ _07570_ _07554_ _07555_ vssd1 vssd1 vccd1 vccd1 _07571_ sky130_fd_sc_hd__mux2_2
XANTENNA__08824__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12764__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10631__B1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17266_ clknet_leaf_133_wb_clk_i _02896_ _00962_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_14478_ net1187 vssd1 vssd1 vccd1 vccd1 _00108_ sky130_fd_sc_hd__inv_2
Xclkload103 clknet_leaf_155_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload103/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_116_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16217_ net1062 vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__inv_2
Xclkload114 clknet_leaf_166_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload114/Y sky130_fd_sc_hd__clkinvlp_4
X_13429_ net2078 net195 net415 vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__mux2_1
Xclkload125 clknet_leaf_171_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload125/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_102_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload136 clknet_leaf_146_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload136/Y sky130_fd_sc_hd__bufinv_16
X_17197_ clknet_leaf_158_wb_clk_i _02827_ _00893_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload147 clknet_leaf_131_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload147/X sky130_fd_sc_hd__clkbuf_8
Xclkload158 clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload158/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_168_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16148_ net1263 vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__inv_2
Xclkload169 clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload169/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_80_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_171_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_171_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13595__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16079_ net1260 vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_100_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08970_ _05026_ _05028_ _05030_ _05032_ vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__or4_1
XANTENNA__09001__B1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08355__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10698__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput1 ACK_I vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12939__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10032__B _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09522_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[3\]
+ net798 net738 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[3\]
+ _05557_ vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__a221o_1
X_09453_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[5\]
+ net852 net843 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05495_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08404_ _04477_ _04479_ _04481_ _04483_ vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09384_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[6\]
+ net611 net606 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__a22o_1
XANTENNA__09068__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08335_ net944 net934 net931 vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__and3_4
XFILLER_0_47_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08815__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout517_A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1259_A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08266_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[25\] _04348_
+ vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__or2_1
X_18333__1322 vssd1 vssd1 vccd1 vccd1 _18333__1322/HI net1322 sky130_fd_sc_hd__conb_1
XFILLER_0_7_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11150__Y _07116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08197_ _04147_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[30\]
+ _04266_ net952 vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__nand4_4
XANTENNA_fanout1047_X net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09240__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout886_A _04281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08594__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1007 net1012 vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__buf_2
X_10090_ _05442_ net365 vssd1 vssd1 vccd1 vccd1 _06118_ sky130_fd_sc_hd__nand2_1
Xfanout1018 net1019 vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__clkbuf_4
Xfanout1029 net1030 vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_10_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout674_X net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09715__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout841_X net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12849__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout939_X net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12800_ net224 net2592 net486 vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__mux2_1
X_13780_ _03749_ _03750_ _03752_ vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__or3_1
XFILLER_0_97_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10992_ _06861_ _06970_ vssd1 vssd1 vccd1 vccd1 _06971_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09846__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12731_ net220 net2282 net495 vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13821__X _03761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15450_ net1149 vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12662_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[27\]
+ net341 vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__and2_1
XFILLER_0_167_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14401_ net1534 vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11613_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[14\] net999 vssd1
+ vssd1 vccd1 vccd1 _07477_ sky130_fd_sc_hd__nand2_2
XFILLER_0_26_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12584__S _03680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15381_ net1080 vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__inv_2
X_12593_ _03612_ net1861 net204 vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17120_ clknet_leaf_129_wb_clk_i _02750_ _00816_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10613__B1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14332_ net375 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11544_ net920 _07418_ _07454_ _07401_ vssd1 vssd1 vccd1 vccd1 _07455_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_137_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17051_ clknet_leaf_191_wb_clk_i _02681_ _00747_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_14263_ _04019_ _04045_ vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__and2b_1
X_11475_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[1\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[1\]
+ net1033 vssd1 vssd1 vccd1 vccd1 _07386_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09609__D net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16002_ net1112 vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__inv_2
X_13214_ net291 net2473 net350 vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__mux2_1
X_10426_ net2527 net258 net540 vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_74_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14194_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[3\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[5\]
+ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[4\] _07027_ vssd1
+ vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__and4_1
XFILLER_0_0_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15196__A net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08585__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13145_ net274 net2747 net446 vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10357_ _06335_ _06376_ net520 vssd1 vssd1 vccd1 vccd1 _06377_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17953_ clknet_leaf_49_wb_clk_i _03292_ _01649_ vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_163_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ net260 net2541 net453 vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_163_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10288_ _06301_ _06303_ _06305_ _06310_ vssd1 vssd1 vccd1 vccd1 _06311_ sky130_fd_sc_hd__or4b_1
X_12027_ _07811_ _07814_ _07832_ _07838_ vssd1 vssd1 vccd1 vccd1 _07839_ sky130_fd_sc_hd__and4bb_1
X_16904_ clknet_leaf_203_wb_clk_i _02534_ _00600_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10133__A _06160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17884_ clknet_leaf_88_wb_clk_i _03227_ _01580_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08742__C1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16835_ clknet_leaf_198_wb_clk_i _02465_ _00531_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12759__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09641__B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13978_ _03848_ _03849_ vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__and2b_1
X_16766_ clknet_leaf_164_wb_clk_i _02396_ _00462_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09298__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09837__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15717_ net1142 vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12929_ _04261_ net562 _03708_ vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__or3_1
X_16697_ clknet_leaf_9_wb_clk_i _02327_ _00393_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_124_Left_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15648_ net1250 vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12494__S _03673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18367_ net1352 vssd1 vssd1 vccd1 vccd1 la_data_out[15] sky130_fd_sc_hd__buf_2
XFILLER_0_8_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15579_ net1249 vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08120_ net1028 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[1\]
+ net972 _04209_ vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__a22o_1
X_17318_ clknet_leaf_115_wb_clk_i _02948_ _01014_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18298_ net1390 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
XFILLER_0_43_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08051_ team_05_WB.instance_to_wrap.total_design.core.data_mem.state\[0\] vssd1 vssd1
+ vccd1 vccd1 _04171_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17249_ clknet_leaf_147_wb_clk_i _02879_ _00945_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09222__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10907__A1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10027__B _06055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08576__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08953_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[15\]
+ net683 net632 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__a22o_1
XANTENNA__08328__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08884_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[17\]
+ net825 net782 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[17\]
+ _04949_ vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__a221o_1
XFILLER_0_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10135__A2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1007_A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout467_A _03710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09289__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09505_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[4\]
+ net641 net612 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout634_A net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08500__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09436_ _05472_ _05474_ _05476_ _05478_ vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__or4_1
XFILLER_0_94_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10702__A1_N team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09367_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[7\]
+ net834 net772 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05413_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout801_A _04394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout422_X net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08318_ _04148_ _04271_ _04365_ net931 vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__and4_4
XFILLER_0_90_842 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12060__A2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09298_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[8\]
+ net667 net658 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05347_ sky130_fd_sc_hd__a22o_1
XANTENNA__09461__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08249_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[31\]
+ net708 net661 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[31\]
+ _04331_ vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__a221o_1
XFILLER_0_144_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12348__B1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11260_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[115\] _07103_
+ _07124_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[27\] vssd1 vssd1
+ vccd1 vccd1 _07222_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_132_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09213__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout791_X net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10211_ _06236_ vssd1 vssd1 vccd1 vccd1 _06237_ sky130_fd_sc_hd__inv_2
XANTENNA__08567__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11191_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[30\] _07124_
+ _07153_ _07155_ vssd1 vssd1 vccd1 vccd1 _07156_ sky130_fd_sc_hd__a211o_1
XANTENNA__10505__X _06518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10374__A2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11571__B2 _07407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10142_ _06166_ _06169_ net514 vssd1 vssd1 vccd1 vccd1 _06170_ sky130_fd_sc_hd__mux2_1
X_10073_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[28\] team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[27\]
+ _06101_ vssd1 vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__and3_1
X_14950_ net1231 vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__inv_2
X_13901_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[22\]
+ net558 net574 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[22\]
+ net985 vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__a221o_1
XANTENNA_input28_A DAT_I[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14881_ net1219 vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__inv_2
XANTENNA__12579__S net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16620_ clknet_leaf_0_wb_clk_i _02250_ _00316_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13832_ net1487 net580 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[10\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__09819__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16551_ clknet_leaf_201_wb_clk_i _02181_ _00247_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13763_ net921 _05921_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[31\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10975_ _06806_ _06807_ _06809_ _06865_ vssd1 vssd1 vccd1 vccd1 _06957_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_69_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15502_ net1172 vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_139_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12714_ net287 net2837 net496 vssd1 vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16482_ clknet_leaf_17_wb_clk_i _02112_ _00178_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13694_ _06771_ _07349_ _03736_ _03735_ _07485_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.next_state\[0\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_57_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18221_ clknet_leaf_79_wb_clk_i net1458 _01916_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_15433_ net1129 vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__inv_2
XANTENNA__13711__B _06572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12645_ team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.state\[1\] team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.state\[0\]
+ net1048 vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_109_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_156_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12587__A0 _03646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13203__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11512__A _07348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15364_ net1227 vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__inv_2
X_18152_ clknet_leaf_19_wb_clk_i _03455_ _01848_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_12576_ _03623_ net1739 net206 vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__mux2_1
XANTENNA__09452__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17103_ clknet_leaf_141_wb_clk_i _02733_ _00799_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_14315_ net377 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[19\]
+ net376 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[18\] vssd1
+ vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__a22oi_2
X_11527_ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[18\] _07437_ net1003
+ vssd1 vssd1 vccd1 vccd1 _07438_ sky130_fd_sc_hd__mux2_2
X_18083_ clknet_leaf_83_wb_clk_i _00010_ _01779_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15295_ net1179 vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14823__A net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17034_ clknet_leaf_17_wb_clk_i _02664_ _00730_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_14246_ _04025_ _04033_ vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__nor2_1
Xhold309 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[105\] vssd1 vssd1
+ vccd1 vccd1 net1723 sky130_fd_sc_hd__dlygate4sd3_1
X_11458_ net919 _07368_ vssd1 vssd1 vccd1 vccd1 _07369_ sky130_fd_sc_hd__nand2_2
XFILLER_0_7_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10409_ _05931_ _05932_ _05973_ vssd1 vssd1 vccd1 vccd1 _06426_ sky130_fd_sc_hd__and3_1
X_14177_ net1936 net503 net909 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[26\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__10562__S net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_4_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11389_ _07315_ _07319_ vssd1 vssd1 vccd1 vccd1 _07320_ sky130_fd_sc_hd__nor2_1
X_13128_ net198 net2133 net445 vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_12__f_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_12__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_13059_ net325 net2799 net456 vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__mux2_1
X_17936_ clknet_leaf_34_wb_clk_i _03275_ _01632_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1009 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2423 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12489__S net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17867_ clknet_leaf_75_wb_clk_i _03210_ _01563_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18332__1321 vssd1 vssd1 vccd1 vccd1 _18332__1321/HI net1321 sky130_fd_sc_hd__conb_1
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_128_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08730__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16818_ clknet_leaf_126_wb_clk_i _02448_ _00514_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_17798_ clknet_leaf_76_wb_clk_i _03141_ _01494_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[108\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_132_Left_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16749_ clknet_leaf_161_wb_clk_i _02379_ _00445_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08555__X team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[26\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09221_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[10\]
+ net771 net751 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[10\]
+ _05272_ vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13113__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09152_ _05203_ _05204_ _05205_ _05206_ vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__or4_1
XANTENNA__12042__A2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[29\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08103_ net1030 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__and2b_1
XANTENNA__14319__A1 _04818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11250__B1 _07120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08797__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12952__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09083_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[13\]
+ net850 net845 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[13\]
+ _05128_ vssd1 vssd1 vccd1 vccd1 _05141_ sky130_fd_sc_hd__a221o_1
XANTENNA__14319__B2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[20\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout215_A _03668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_141_Left_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08034_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[15\] vssd1
+ vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__inv_2
Xinput70 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold810 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2224 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold821 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net2235 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold832 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net2246 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold843 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 net2257 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08549__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold854 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2268 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold865 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 net2279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold898 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2312 sky130_fd_sc_hd__dlygate4sd3_1
X_09985_ net373 net361 vssd1 vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08936_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[16\]
+ net794 net733 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__a22o_1
Xhold1510 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 net2924 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1521 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 net2935 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12399__S _07852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1532 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 net2946 sky130_fd_sc_hd__dlygate4sd3_1
X_08867_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[17\]
+ net703 net640 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[17\]
+ _04926_ vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__a221o_1
Xhold1543 team_05_WB.instance_to_wrap.total_design.keypad0.key_counter\[0\] vssd1
+ vssd1 vccd1 vccd1 net2957 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout372_X net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_150_Left_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1554 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net2968 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout849_A _04370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08721__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08798_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[19\]
+ net844 net733 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09712__D net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09512__A_N net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_8_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout637_X net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10760_ net334 _06324_ _06755_ _06757_ vssd1 vssd1 vccd1 vccd1 _06758_ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09419_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[6\]
+ net590 _05462_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[6\]
+ sky130_fd_sc_hd__o21a_4
XFILLER_0_66_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10691_ _06413_ net347 vssd1 vssd1 vccd1 vccd1 _06693_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_203_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_203_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout804_X net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13023__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12430_ _03665_ net1854 _03668_ vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__mux2_1
XANTENNA__14346__C _04094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09434__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11241__B1 _07109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12361_ _07884_ _08022_ _03549_ _03603_ vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__o22a_1
XFILLER_0_117_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12862__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14100_ _03956_ _03965_ vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11312_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[48\] _07117_
+ _07121_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[80\] vssd1 vssd1
+ vccd1 vccd1 _07271_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15080_ net1224 vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__inv_2
XANTENNA__09737__A _05768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12292_ _03579_ _03582_ _03578_ vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__o21ai_1
X_14031_ _03866_ _03871_ _03900_ vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11243_ _07201_ _07203_ _07204_ _07205_ vssd1 vssd1 vccd1 vccd1 _07206_ sky130_fd_sc_hd__or4_1
XANTENNA__11544__A1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11174_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[15\] _07101_
+ _07130_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[103\] _07139_
+ vssd1 vssd1 vccd1 vccd1 _07140_ sky130_fd_sc_hd__a221o_1
XANTENNA__08960__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10125_ net377 net364 vssd1 vssd1 vccd1 vccd1 _06153_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15982_ net1140 vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__inv_2
X_17721_ clknet_leaf_100_wb_clk_i _03064_ _01417_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[95\]
+ sky130_fd_sc_hd__dfrtp_1
X_10056_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[3\] team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06085_ sky130_fd_sc_hd__nand2_1
X_14933_ net1079 vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18407__1375 vssd1 vssd1 vccd1 vccd1 _18407__1375/HI net1375 sky130_fd_sc_hd__conb_1
XANTENNA__08712__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17652_ clknet_leaf_39_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[19\]
+ _01348_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_14864_ net1093 vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16603_ clknet_leaf_193_wb_clk_i _02233_ _00299_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13815_ net1676 net969 net723 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[26\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_159_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17583_ clknet_leaf_73_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[20\]
+ _01279_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_14795_ net1067 vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_158_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13722__A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13746_ _05213_ _06521_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[14\]
+ sky130_fd_sc_hd__nor2_1
X_16534_ clknet_leaf_139_wb_clk_i _02164_ _00230_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10958_ _06943_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[20\] net564
+ vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16465_ clknet_leaf_169_wb_clk_i _02095_ _00161_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13677_ net2446 net284 net384 vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__mux2_1
X_10889_ _06778_ _06885_ _06775_ _06776_ vssd1 vssd1 vccd1 vccd1 _06886_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_85_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18204_ clknet_leaf_36_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[25\]
+ _01899_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12628_ _03632_ net1811 net201 vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15416_ net1113 vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16396_ clknet_leaf_2_wb_clk_i _02026_ _00092_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09425__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11232__B1 _07097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15347_ net1213 vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__inv_2
XANTENNA__08779__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18135_ clknet_leaf_32_wb_clk_i _03438_ _01831_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_171_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12559_ _03612_ net1835 net205 vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__mux2_1
XANTENNA__12772__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18066_ clknet_leaf_86_wb_clk_i _03404_ _01762_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__dfrtp_1
Xhold106 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[27\]
+ vssd1 vssd1 vccd1 vccd1 net1520 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15278_ net1190 vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__inv_2
Xhold117 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[5\] vssd1 vssd1
+ vccd1 vccd1 net1531 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold128 team_05_WB.instance_to_wrap.total_design.key_data vssd1 vssd1 vccd1 vccd1
+ net1542 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14229_ team_05_WB.instance_to_wrap.total_design.keypad0.counter\[13\] team_05_WB.instance_to_wrap.total_design.keypad0.counter\[14\]
+ _04024_ vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__and3_1
Xhold139 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[15\]
+ vssd1 vssd1 vccd1 vccd1 net1553 sky130_fd_sc_hd__dlygate4sd3_1
X_17017_ clknet_leaf_6_wb_clk_i _02647_ _00713_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_78_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08270__B team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[20\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout608 _04320_ vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout619 net620 vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__buf_4
XANTENNA__15384__A net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12360__X _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09770_ _05795_ _05797_ _05800_ net716 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__o32a_2
XFILLER_0_77_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08721_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[22\]
+ net800 net791 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__a22o_1
XANTENNA__11299__B1 _07121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17919_ clknet_leaf_40_wb_clk_i _03258_ _01615_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.BUSY_O
+ sky130_fd_sc_hd__dfrtp_2
Xfanout1190 net1211 vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__buf_2
XANTENNA__13108__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08652_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[23\]
+ net618 net616 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[23\]
+ _04719_ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__a221o_1
XFILLER_0_135_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10510__A2 _06521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08583_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[25\]
+ net823 net757 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__a22o_1
XANTENNA__12947__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08285__X _04367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08726__A _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09204_ net953 _04352_ _04269_ vssd1 vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__a21o_1
XANTENNA__14166__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09416__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11223__B1 _07121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09135_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[11\]
+ net703 net699 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1241_A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09066_ _04354_ _05124_ vssd1 vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout799_A net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold640 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 net2054 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold651 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net2065 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1127_X net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09707__D net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold662 net133 vssd1 vssd1 vccd1 vccd1 net2076 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold673 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2087 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09195__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold684 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[116\] vssd1 vssd1
+ vccd1 vccd1 net2098 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold695 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net2109 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15294__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09563__Y team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09968_ _05914_ _05927_ vssd1 vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__or2_1
X_08919_ _04977_ _04979_ _04981_ _04983_ vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__or4_1
XANTENNA_clkbuf_leaf_83_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09899_ _04613_ _04632_ vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout754_X net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09723__C net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1340 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2754 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13018__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11930_ _07698_ _07707_ vssd1 vssd1 vccd1 vccd1 _07742_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_86_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1351 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2765 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1362 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2776 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1373 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2787 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1384 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2798 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1395 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 net2809 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08339__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout921_X net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11861_ _07636_ _07648_ vssd1 vssd1 vccd1 vccd1 _07673_ sky130_fd_sc_hd__xnor2_2
XANTENNA__12857__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14638__A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13600_ net1996 net234 net394 vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10812_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[15\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06809_ sky130_fd_sc_hd__and2_1
XFILLER_0_170_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14580_ net1068 vssd1 vssd1 vccd1 vccd1 _00210_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09655__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11792_ _07603_ vssd1 vssd1 vccd1 vccd1 _07604_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_101_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13531_ net1981 net224 net402 vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10743_ _05735_ _05944_ vssd1 vssd1 vccd1 vccd1 _06742_ sky130_fd_sc_hd__xor2_1
XFILLER_0_137_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16250_ net1138 vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13462_ net196 net2087 net410 vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__mux2_1
X_10674_ _05507_ net552 _06676_ vssd1 vssd1 vccd1 vccd1 _06677_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_11_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09407__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15201_ net1228 vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__inv_2
X_12413_ net1712 _07793_ _03667_ vssd1 vssd1 vccd1 vccd1 _03217_ sky130_fd_sc_hd__mux2_1
XANTENNA__11214__B1 _07127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13688__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16181_ net1134 vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__inv_2
XANTENNA__12592__S net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13393_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[0\]
+ net305 net423 vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__mux2_1
X_18331__1320 vssd1 vssd1 vccd1 vccd1 _18331__1320/HI net1320 sky130_fd_sc_hd__conb_1
X_15132_ net1095 vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12344_ _07774_ net354 _03530_ _03540_ vssd1 vssd1 vccd1 vccd1 _03639_ sky130_fd_sc_hd__o31a_1
XFILLER_0_121_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15063_ net1101 vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12275_ _03564_ _03566_ _07978_ vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09617__D net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14014_ net979 net980 vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__nand2b_1
X_11226_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[124\] _07099_
+ _07126_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[84\] vssd1 vssd1
+ vccd1 vccd1 _07189_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09186__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08394__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13717__A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08933__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11157_ _07039_ _07122_ vssd1 vssd1 vccd1 vccd1 _07123_ sky130_fd_sc_hd__nor2_4
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09914__B net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_147_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10108_ _05165_ net365 vssd1 vssd1 vccd1 vccd1 _06136_ sky130_fd_sc_hd__nand2_1
X_11088_ _07043_ _07054_ _07048_ vssd1 vssd1 vccd1 vccd1 _07055_ sky130_fd_sc_hd__o21ai_1
X_15965_ net1269 vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__inv_2
X_17704_ clknet_leaf_93_wb_clk_i _03047_ _01400_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[78\]
+ sky130_fd_sc_hd__dfrtp_1
X_14916_ net1235 vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__inv_2
X_10039_ _04533_ net363 vssd1 vssd1 vccd1 vccd1 _06068_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_125_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_196_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_196_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15896_ net1266 vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13690__A1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17635_ clknet_leaf_70_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[2\]
+ _01331_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14847_ net1178 vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__inv_2
XANTENNA__12767__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_125_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_125_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_19_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13442__A1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17566_ clknet_leaf_113_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[3\]
+ _01262_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_14778_ net1055 vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09110__A2 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16517_ clknet_leaf_176_wb_clk_i _02147_ _00213_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_173_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13729_ net899 _06185_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[29\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17497_ clknet_leaf_114_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[0\]
+ _01193_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_129_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08265__B net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_128_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16448_ clknet_leaf_131_wb_clk_i _02078_ _00144_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_144_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09088__A_N _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13598__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14283__A _06540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12355__X _03650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16379_ clknet_leaf_191_wb_clk_i _02009_ _00075_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18118_ clknet_leaf_46_wb_clk_i _00032_ _01814_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18049_ net1039 _03387_ _01745_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09177__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10035__B net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout405 net406 vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_39_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout416 _03726_ vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__buf_6
X_09822_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[20\]
+ net617 net614 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[20\]
+ _05842_ vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__a221o_1
Xfanout427 _03724_ vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__buf_4
XANTENNA__08924__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout438 _03721_ vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__buf_6
Xfanout449 _03714_ vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__buf_4
X_09753_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[0\]
+ net887 net866 _04296_ vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_33_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08704_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[22\]
+ net718 _04770_ _04776_ vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_146_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09684_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[1\]
+ net883 net867 net860 vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__and4_1
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08635_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[24\]
+ net796 net734 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[24\]
+ _04699_ vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_167_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_96_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08566_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[25\]
+ net638 net631 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11153__Y _07119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09101__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08497_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[27\]
+ net803 net788 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout714_A _04288_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1012 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13197__A0 _06247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14193__A _07031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1244_X net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13301__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09118_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[12\]
+ net813 net733 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__a22o_1
X_10390_ _05841_ _05884_ vssd1 vssd1 vccd1 vccd1 _06408_ sky130_fd_sc_hd__xnor2_4
XANTENNA__08191__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[14\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09718__C net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09049_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[13\]
+ net668 net629 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__a22o_1
XANTENNA__14921__A net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09168__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12060_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[11\] team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[13\]
+ net998 net543 vssd1 vssd1 vccd1 vccd1 _07872_ sky130_fd_sc_hd__a31oi_1
Xhold470 team_05_WB.instance_to_wrap.total_design.core.data_mem.state\[2\] vssd1 vssd1
+ vccd1 vccd1 net1884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[35\] vssd1 vssd1
+ vccd1 vccd1 net1895 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout871_X net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17654__D team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[21\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08376__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11011_ _06986_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[10\] net568
+ vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__mux2_1
Xhold492 team_05_WB.instance_to_wrap.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 net1906
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11609__X _07475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08915__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10513__X _06525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout950 _04363_ vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__buf_2
Xfanout961 net962 vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__clkbuf_4
Xfanout972 net973 vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__buf_1
Xfanout983 net984 vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__buf_2
Xfanout994 _07470_ vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15750_ net1272 vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__inv_2
X_12962_ net563 _03695_ _03708_ vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__or3_4
Xhold1170 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2584 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input10_A DAT_I[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09340__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14701_ net1082 vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__inv_2
Xhold1181 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net2595 sky130_fd_sc_hd__dlygate4sd3_1
X_11913_ _07702_ _07705_ vssd1 vssd1 vccd1 vccd1 _07725_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_142_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1192 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2606 sky130_fd_sc_hd__dlygate4sd3_1
X_15681_ net1149 vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__inv_2
XANTENNA__12587__S _03681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12893_ net308 net2772 net479 vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17420_ clknet_leaf_50_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[20\]
+ _01116_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14632_ net1224 vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ _07623_ _07628_ vssd1 vssd1 vccd1 vccd1 _07656_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09628__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17351_ clknet_leaf_37_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[15\]
+ _01047_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_14563_ net1204 vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__inv_2
X_11775_ _07449_ _07523_ vssd1 vssd1 vccd1 vccd1 _07587_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16302_ net1155 vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13514_ net2274 net292 net404 vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__mux2_1
X_10726_ _06663_ _06725_ net527 vssd1 vssd1 vccd1 vccd1 _06726_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14494_ net1062 vssd1 vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__inv_2
X_17282_ clknet_leaf_6_wb_clk_i _02912_ _00978_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_16233_ net1136 vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13445_ net2149 net274 net414 vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10657_ _06118_ _06130_ vssd1 vssd1 vccd1 vccd1 _06661_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13211__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload15 clknet_leaf_200_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload15/Y sky130_fd_sc_hd__inv_6
XFILLER_0_35_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload26 clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload26/Y sky130_fd_sc_hd__clkinv_2
X_16164_ net1152 vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__inv_2
Xclkload37 clknet_leaf_186_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload37/Y sky130_fd_sc_hd__clkinvlp_4
X_13376_ net2255 net259 net423 vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_118_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10588_ _06524_ _06595_ net529 vssd1 vssd1 vccd1 vccd1 _06596_ sky130_fd_sc_hd__mux2_1
XANTENNA__10407__Y _06424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload48 clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload48/Y sky130_fd_sc_hd__bufinv_16
Xclkload59 clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload59/Y sky130_fd_sc_hd__clkinv_16
X_12327_ _03531_ _03540_ net543 vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__a21oi_2
X_15115_ net1076 vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_77_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16095_ net1307 vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__inv_2
XANTENNA__10136__A _04613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09159__A2 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15046_ net1209 vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__inv_2
XFILLER_0_167_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12258_ _07880_ _07891_ _07871_ vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__a21boi_1
XANTENNA__08367__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17564__D team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11209_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[77\] _07109_
+ _07128_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[69\] _07172_
+ vssd1 vssd1 vccd1 vccd1 _07173_ sky130_fd_sc_hd__a221o_1
XANTENNA__08906__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09644__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12189_ _07941_ _07986_ _07981_ vssd1 vssd1 vccd1 vccd1 _08001_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_166_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10713__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16997_ clknet_leaf_180_wb_clk_i _02627_ _00693_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_15948_ net1303 vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__inv_2
XANTENNA__12497__S _03673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15879_ net1292 vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__inv_2
X_08420_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[29\]
+ net850 net785 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[29\]
+ _04496_ vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__a221o_1
X_17618_ clknet_leaf_58_wb_clk_i _02989_ _01314_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08351_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[30\]
+ net677 net626 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[30\]
+ _04431_ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__a221o_1
X_17549_ clknet_leaf_58_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[20\]
+ _01245_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08282_ _04237_ _04241_ _04148_ _04231_ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__a211o_1
Xclkload9 clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload9/Y sky130_fd_sc_hd__inv_8
XFILLER_0_73_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_93_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12926__A0 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13121__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_22_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08070__A2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[26\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12960__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10046__A _04613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10952__A2 _06387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08358__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout202 _03683_ vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__buf_4
XANTENNA_fanout497_A net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout213 _03671_ vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__buf_4
Xfanout224 net225 vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__buf_2
Xfanout235 net237 vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__clkbuf_2
Xfanout246 net249 vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input2_A DAT_I[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09805_ _05104_ _05834_ _05057_ _05102_ vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__a211o_1
Xfanout257 _06442_ vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_31_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout268 _06499_ vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout279 net281 vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout664_A _04305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09736_ _05764_ _05766_ _05767_ _05737_ vssd1 vssd1 vccd1 vccd1 _05768_ sky130_fd_sc_hd__a31o_2
XFILLER_0_69_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09322__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09667_ net572 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[1\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[1\] vssd1 vssd1 vccd1
+ vccd1 _05700_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout452_X net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout831_A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11164__X _07130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08530__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_19_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08618_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[24\]
+ net608 _04692_ net721 vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__a211o_1
XFILLER_0_55_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09598_ net571 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[2\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[2\] vssd1 vssd1 vccd1
+ vccd1 _05633_ sky130_fd_sc_hd__a21oi_2
XANTENNA__09720__D net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08549_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[26\]
+ net812 net753 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[26\]
+ _04625_ vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout717_X net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11560_ net1778 net1004 _07441_ net358 vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08294__C1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[20\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17649__D team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[16\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10511_ net518 _06133_ _06146_ vssd1 vssd1 vccd1 vccd1 _06523_ sky130_fd_sc_hd__and3_1
XFILLER_0_134_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11491_ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[22\] _07400_ net1001
+ vssd1 vssd1 vccd1 vccd1 _07402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08192__Y _04275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13031__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13230_ net199 net2740 net439 vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__mux2_1
X_10442_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[18\] _06095_ vssd1
+ vssd1 vccd1 vccd1 _06458_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09389__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11196__A2 _07125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12393__A1 _03605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08597__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13161_ net200 net2630 net442 vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__mux2_1
X_10373_ _04839_ _06391_ vssd1 vssd1 vccd1 vccd1 _06392_ sky130_fd_sc_hd__nand2_1
XANTENNA__12870__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12112_ _07923_ vssd1 vssd1 vccd1 vccd1 _07924_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input58_A wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13092_ net326 net1984 net453 vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08349__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11486__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12043_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[23\] team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[25\]
+ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[26\] team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[28\]
+ net993 vssd1 vssd1 vccd1 vccd1 _07855_ sky130_fd_sc_hd__o41a_1
X_16920_ clknet_leaf_27_wb_clk_i _02550_ _00616_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16851_ clknet_leaf_164_wb_clk_i _02481_ _00547_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout780 net781 vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__buf_4
X_15802_ net1298 vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__inv_2
Xfanout791 net793 vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_4_14__f_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16782_ clknet_leaf_178_wb_clk_i _02412_ _00478_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_161_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13994_ _03863_ _03864_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__nand2_1
XANTENNA__09849__B1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[21\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_161_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10459__A1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09313__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15733_ net1269 vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__inv_2
XANTENNA__10459__B2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13714__B _06521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12945_ net267 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[16\]
+ net468 vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08521__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13206__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15664_ net1155 vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12876_ net260 net2220 net479 vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__mux2_1
X_17403_ clknet_leaf_56_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[3\]
+ _01099_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10776__D team_05_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14615_ net1101 vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18383_ net1368 vssd1 vssd1 vccd1 vccd1 la_data_out[31] sky130_fd_sc_hd__buf_2
X_11827_ _07615_ _07617_ _07638_ _07590_ vssd1 vssd1 vccd1 vccd1 _07639_ sky130_fd_sc_hd__a31o_1
X_15595_ net1161 vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13730__A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17334_ clknet_leaf_140_wb_clk_i _02964_ _01030_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11758_ _07554_ _07557_ vssd1 vssd1 vccd1 vccd1 _07570_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14546_ net1238 vssd1 vssd1 vccd1 vccd1 _00176_ sky130_fd_sc_hd__inv_2
XANTENNA__08285__C1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10631__A1 _04174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10709_ net516 _06678_ vssd1 vssd1 vccd1 vccd1 _06710_ sky130_fd_sc_hd__nor2_1
X_17265_ clknet_leaf_169_wb_clk_i _02895_ _00961_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11689_ net63 net62 _07501_ _07502_ vssd1 vssd1 vccd1 vccd1 _07503_ sky130_fd_sc_hd__or4_1
X_14477_ net1087 vssd1 vssd1 vccd1 vccd1 _00107_ sky130_fd_sc_hd__inv_2
XANTENNA__09639__B net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload104 clknet_leaf_156_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload104/X sky130_fd_sc_hd__clkbuf_8
X_16216_ net1057 vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13428_ net2160 net198 net415 vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__mux2_1
Xclkload115 clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload115/X sky130_fd_sc_hd__clkbuf_4
X_17196_ clknet_leaf_7_wb_clk_i _02826_ _00892_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload126 clknet_leaf_172_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload126/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_12_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload137 clknet_leaf_147_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload137/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__11187__A2 _07102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12384__A1 _03645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload148 clknet_leaf_133_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload148/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__08588__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload159 clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload159/Y sky130_fd_sc_hd__inv_6
X_16147_ net1263 vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_168_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10395__A0 _06237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12780__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13359_ net325 net2929 net425 vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_168_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16078_ net1260 vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15029_ net1060 vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10698__A1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09552__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_140_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_140_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08760__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput2 DAT_I[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09521_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[3\]
+ net760 net756 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08512__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13116__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09452_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[5\]
+ net808 net753 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05494_ sky130_fd_sc_hd__a22o_1
XANTENNA__11426__B1_N net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08403_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[29\]
+ net703 net681 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[29\]
+ _04482_ vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09383_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[6\]
+ net618 net602 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__a22o_1
XANTENNA__12955__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout245_A _06294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08334_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[31\]
+ net753 net749 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[31\]
+ _04413_ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__a221o_1
XFILLER_0_52_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08293__X _04375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10083__C1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08265_ _04148_ net1017 vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_864 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout412_A _03727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08196_ _04147_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[30\]
+ _04266_ _04278_ vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__and4_2
XANTENNA__12375__A1 _07793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11178__A2 _07091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12543__X _03678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_93_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_93_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout879_A net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1008 net1009 vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__buf_2
Xfanout1019 net1021 vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__buf_2
XANTENNA__09715__D net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09543__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout667_X net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08751__B1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08643__A_N net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_27_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09719_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[0\]
+ net1017 net951 net934 vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__and4_1
X_10991_ _06813_ _06815_ vssd1 vssd1 vccd1 vccd1 _06970_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout834_X net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08503__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13026__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12730_ net190 net2540 net495 vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__mux2_1
XANTENNA__10310__B1 _06055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12661_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[28\]
+ net342 vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__and2_1
XANTENNA__12865__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14400_ net1507 vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11612_ net1603 net1009 _07472_ _07476_ vssd1 vssd1 vccd1 vccd1 _03308_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12592_ _03614_ net1893 net204 vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__mux2_1
X_15380_ net1075 vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11543_ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[22\] net1001 _07349_
+ _07351_ team_05_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 _07454_ sky130_fd_sc_hd__o221a_1
XFILLER_0_25_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14331_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[1\] _05732_
+ vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_137_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_36_Left_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14262_ team_05_WB.instance_to_wrap.total_design.keypad0.counter\[3\] team_05_WB.instance_to_wrap.total_design.keypad0.counter\[4\]
+ _04017_ team_05_WB.instance_to_wrap.total_design.keypad0.counter\[5\] vssd1 vssd1
+ vccd1 vccd1 _04045_ sky130_fd_sc_hd__a31o_1
X_17050_ clknet_leaf_31_wb_clk_i _02680_ _00746_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11474_ net1050 net1049 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[1\]
+ vssd1 vssd1 vccd1 vccd1 _07385_ sky130_fd_sc_hd__o21a_1
XFILLER_0_107_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11169__A2 _07113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12366__A1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13213_ _06570_ net2655 net350 vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__mux2_1
X_16001_ net1112 vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10425_ _06437_ _06441_ net382 vssd1 vssd1 vccd1 vccd1 _06442_ sky130_fd_sc_hd__o21a_4
X_14193_ _07031_ net729 _03999_ vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_74_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13144_ net270 net2882 net444 vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10356_ _06149_ _06168_ vssd1 vssd1 vccd1 vccd1 _06376_ sky130_fd_sc_hd__nand2_1
XANTENNA__13709__B _06609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17465__Q team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_11__f_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_11__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__08990__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17952_ clknet_leaf_52_wb_clk_i net2819 _01648_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__dfrtp_1
X_13075_ net265 net2930 net452 vssd1 vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__mux2_1
X_10287_ net336 _06308_ _06309_ net337 vssd1 vssd1 vccd1 vccd1 _06310_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_163_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14287__D_N _06320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12026_ _07834_ _07835_ _07837_ _07799_ vssd1 vssd1 vccd1 vccd1 _07838_ sky130_fd_sc_hd__o22a_1
X_16903_ clknet_leaf_203_wb_clk_i _02533_ _00599_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09534__A2 _04366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17883_ clknet_leaf_75_wb_clk_i _03226_ _01579_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08742__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_45_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16834_ clknet_leaf_8_wb_clk_i _02464_ _00530_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16765_ clknet_leaf_108_wb_clk_i _02395_ _00461_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13977_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[9\] _03824_ _03823_
+ vssd1 vssd1 vccd1 vccd1 _03849_ sky130_fd_sc_hd__a21bo_1
XANTENNA__09641__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15716_ net1142 vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__inv_2
X_12928_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[9\] _04254_
+ vssd1 vssd1 vccd1 vccd1 _03708_ sky130_fd_sc_hd__or2_2
XFILLER_0_158_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16696_ clknet_leaf_33_wb_clk_i _02326_ _00392_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10852__A1 _06847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15647_ net1243 vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__inv_2
XANTENNA__12775__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12859_ net324 net2810 net483 vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13460__A team_05_WB.instance_to_wrap.total_design.core.instr_fetch vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18366_ net1351 vssd1 vssd1 vccd1 vccd1 la_data_out[14] sky130_fd_sc_hd__buf_2
X_15578_ net1249 vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17317_ clknet_leaf_176_wb_clk_i _02947_ _01013_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[13\]
+ sky130_fd_sc_hd__dfrtp_2
X_14529_ net1236 vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__inv_2
X_18297_ net1389 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
XANTENNA__09470__B2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[11\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08050_ net1648 vssd1 vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17248_ clknet_leaf_131_wb_clk_i _02878_ _00944_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17179_ clknet_leaf_193_wb_clk_i _02809_ _00875_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14291__A _04573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10907__A2 _06185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08981__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08952_ _05014_ vssd1 vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__inv_2
XANTENNA__09525__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08883_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[17\]
+ net787 net768 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09911__A_N net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08733__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08288__X _04370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout362_A _05770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09504_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[4\]
+ net692 net595 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[4\]
+ _05542_ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_13__f_wb_clk_i_X clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_17_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09435_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[5\]
+ net709 net631 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[5\]
+ _05477_ vssd1 vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1271_A net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout627_A net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09366_ _05405_ _05407_ _05409_ _05411_ vssd1 vssd1 vccd1 vccd1 _05412_ sky130_fd_sc_hd__or4_1
XFILLER_0_164_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13801__C net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12596__A1 _07812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11161__Y _07127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08317_ _04379_ _04386_ _04392_ _04398_ vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_43_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09297_ _05339_ _05341_ _05343_ _05345_ vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout415_X net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08248_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[31\]
+ net666 net642 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout996_A _07470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15297__A net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08179_ _04254_ _04255_ vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_132_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10210_ _05634_ _06235_ vssd1 vssd1 vccd1 vccd1 _06236_ sky130_fd_sc_hd__nor2_1
XFILLER_0_162_1068 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11020__A1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11190_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[46\] _07091_
+ _07100_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[6\] _07154_
+ vssd1 vssd1 vccd1 vccd1 _07155_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_1154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout784_X net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10241__A1_N _06049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10141_ _06167_ _06168_ vssd1 vssd1 vccd1 vccd1 _06169_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput180 net180 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__clkbuf_4
XANTENNA__18401__A net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10072_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[26\] _06100_ vssd1
+ vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout951_X net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11323__A2 _07115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12520__A1 _03610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13900_ net1548 net981 _03786_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[21\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__08198__X _04281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14880_ net1105 vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13831_ net1465 net582 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[9\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_173_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16550_ clknet_leaf_118_wb_clk_i _02180_ _00246_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13762_ net921 _06108_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[30\]
+ sky130_fd_sc_hd__nor2_1
X_10974_ _06956_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[17\] net564
+ vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15501_ net1164 vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_139_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12713_ net290 net2950 net496 vssd1 vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__mux2_1
XANTENNA__12595__S _03681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16481_ clknet_leaf_151_wb_clk_i _02111_ _00177_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13693_ team_05_WB.EN_VAL_REG _00040_ net1048 team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_139_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18220_ clknet_leaf_80_wb_clk_i net1585 _01915_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_15432_ net1115 vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__inv_2
X_12644_ _03623_ net1788 net201 vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_156_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_156_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18151_ clknet_leaf_196_wb_clk_i _03454_ _01847_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12575_ _03641_ net1806 net205 vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__mux2_1
X_15363_ net1197 vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08255__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17102_ clknet_leaf_169_wb_clk_i _02732_ _00798_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14314_ net360 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[20\]
+ vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__nor2_1
X_11526_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[18\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[18\]
+ net1031 vssd1 vssd1 vccd1 vccd1 _07437_ sky130_fd_sc_hd__mux2_1
X_18082_ clknet_leaf_83_wb_clk_i _00009_ _01778_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_15294_ net1063 vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17033_ clknet_leaf_21_wb_clk_i _02663_ _00729_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14245_ team_05_WB.instance_to_wrap.total_design.keypad0.counter\[13\] _04024_ net2526
+ vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__a21oi_1
X_11457_ net920 _07365_ vssd1 vssd1 vccd1 vccd1 _07368_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10408_ net889 _06424_ vssd1 vssd1 vccd1 vccd1 _06425_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14176_ net1725 net503 net908 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[25\]
+ sky130_fd_sc_hd__and3_1
X_11388_ _07312_ _07316_ _07317_ _07318_ vssd1 vssd1 vccd1 vccd1 _07319_ sky130_fd_sc_hd__or4_1
XANTENNA__08963__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15935__A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10339_ _06060_ _06359_ net372 vssd1 vssd1 vccd1 vccd1 _06360_ sky130_fd_sc_hd__mux2_1
X_13127_ _04257_ net562 _03698_ vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__or3_1
X_17935_ clknet_leaf_34_wb_clk_i _03274_ _01631_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13058_ net322 net2847 net456 vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_9__f_wb_clk_i_X clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12511__A1 _03661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11314__A2 _07092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08715__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17572__D team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11527__X _07438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12009_ _07516_ _07623_ _07820_ vssd1 vssd1 vccd1 vccd1 _07821_ sky130_fd_sc_hd__o21a_2
X_17866_ clknet_leaf_98_wb_clk_i _03209_ _01562_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09652__B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16817_ clknet_leaf_172_wb_clk_i _02447_ _00513_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17797_ clknet_leaf_103_wb_clk_i _03140_ _01493_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[107\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08268__B team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[27\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_34_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16748_ clknet_leaf_4_wb_clk_i _02378_ _00444_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09140__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14286__A _06369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16679_ clknet_leaf_202_wb_clk_i _02309_ _00375_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09220_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[10\]
+ net756 net741 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09151_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[11\]
+ net691 net621 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[11\]
+ _05190_ vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18349_ net1334 vssd1 vssd1 vccd1 vccd1 irq[0] sky130_fd_sc_hd__buf_2
XFILLER_0_17_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08246__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12042__A3 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[30\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10589__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08102_ net1029 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[10\]
+ net974 _04200_ vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09082_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[13\]
+ net774 net736 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[13\]
+ _05130_ vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__a221o_1
XANTENNA__14319__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[21\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10053__A2 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10038__B _05770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14341__A2_N net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08033_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[16\] vssd1
+ vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput60 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__buf_1
Xhold800 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2214 sky130_fd_sc_hd__dlygate4sd3_1
Xinput71 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold811 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2225 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout208_A _03676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold822 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2236 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold833 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net2258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold855 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2280 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08954__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold877 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2291 sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 net2302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold899 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2313 sky130_fd_sc_hd__dlygate4sd3_1
X_09984_ net374 net366 vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08935_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[16\]
+ net756 net745 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[16\]
+ _04998_ vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_73_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12502__A1 _07821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1500 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2914 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08706__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1511 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net2925 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1522 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[6\] vssd1 vssd1
+ vccd1 vccd1 net2936 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1533 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 net2947 sky130_fd_sc_hd__dlygate4sd3_1
X_08866_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[17\]
+ net691 net621 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[17\]
+ _04932_ vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__a221o_1
Xhold1544 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2958 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1555 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2969 sky130_fd_sc_hd__dlygate4sd3_1
X_08797_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[19\]
+ net827 net763 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[19\]
+ _04862_ vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_88_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11608__A3 _07472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout911_A net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08485__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11613__A team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[14\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13304__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09418_ _05448_ _05449_ _05457_ _05461_ vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__or4_1
X_10690_ net890 _06691_ _06690_ net555 vssd1 vssd1 vccd1 vccd1 _06692_ sky130_fd_sc_hd__a211o_1
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08194__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[27\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09349_ _05381_ _05382_ _05394_ _05395_ vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_134_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12360_ net354 _03608_ _03616_ _07474_ vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__o22a_2
XFILLER_0_105_411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11311_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[24\] _07119_
+ _07120_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[32\] _07269_
+ vssd1 vssd1 vccd1 vccd1 _07270_ sky130_fd_sc_hd__a221o_1
XANTENNA__10638__A2_N _06051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12291_ _03512_ _03585_ vssd1 vssd1 vccd1 vccd1 _03586_ sky130_fd_sc_hd__nor2_1
X_14030_ _03898_ _03899_ vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__nand2b_1
XANTENNA__09198__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11242_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[4\] _07100_ _07105_
+ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[12\] _07195_ vssd1 vssd1
+ vccd1 vccd1 _07205_ sky130_fd_sc_hd__a221o_1
XANTENNA__08945__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11173_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[23\] _07125_
+ _07129_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[63\] vssd1 vssd1
+ vccd1 vccd1 _07139_ sky130_fd_sc_hd__a22o_1
XANTENNA__10752__B1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input40_A wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10124_ net367 net360 vssd1 vssd1 vccd1 vccd1 _06152_ sky130_fd_sc_hd__nand2_1
X_15981_ net1173 vssd1 vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17720_ clknet_leaf_93_wb_clk_i _03063_ _01416_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[94\]
+ sky130_fd_sc_hd__dfrtp_1
X_10055_ _06001_ _06083_ _04275_ vssd1 vssd1 vccd1 vccd1 _06084_ sky130_fd_sc_hd__o21a_1
X_14932_ net1069 vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__inv_2
XANTENNA__09370__B1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17651_ clknet_leaf_39_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[18\]
+ _01347_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_14863_ net1280 vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16602_ clknet_leaf_11_wb_clk_i _02232_ _00298_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13814_ net1667 net969 net723 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[25\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_98_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17582_ clknet_leaf_73_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[19\]
+ _01278_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_14794_ net1122 vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_158_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09122__B1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16533_ clknet_leaf_23_wb_clk_i _02163_ _00229_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13745_ net922 _06540_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[13\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__13722__B _06369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10957_ net956 _06408_ _06942_ vssd1 vssd1 vccd1 vccd1 _06943_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_123_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13214__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16464_ clknet_leaf_138_wb_clk_i _02094_ _00160_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_118_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13676_ net2342 net275 net386 vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__mux2_1
X_10888_ _06777_ _06884_ vssd1 vssd1 vccd1 vccd1 _06885_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18203_ clknet_leaf_35_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[24\]
+ _01898_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_15415_ net1131 vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12627_ _03612_ net1839 net202 vssd1 vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16395_ clknet_leaf_187_wb_clk_i _02025_ _00091_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10139__A net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18134_ clknet_leaf_47_wb_clk_i _00030_ _01830_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_171_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15346_ net1232 vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12558_ _03614_ net1793 net205 vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_171_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17567__D team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18065_ clknet_leaf_86_wb_clk_i _03403_ _01761_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__dfrtp_1
X_11509_ _07399_ _07410_ _07419_ vssd1 vssd1 vccd1 vccd1 _07420_ sky130_fd_sc_hd__or3_1
XFILLER_0_124_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15277_ net1081 vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09647__B net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold107 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[20\]
+ vssd1 vssd1 vccd1 vccd1 net1521 sky130_fd_sc_hd__dlygate4sd3_1
X_12489_ net1684 _03614_ net211 vssd1 vssd1 vccd1 vccd1 _03147_ sky130_fd_sc_hd__mux2_1
Xhold118 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[0\]
+ vssd1 vssd1 vccd1 vccd1 net1532 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09189__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17016_ clknet_leaf_29_wb_clk_i _02646_ _00712_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold129 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1543 sky130_fd_sc_hd__dlygate4sd3_1
X_14228_ team_05_WB.instance_to_wrap.total_design.keypad0.counter\[12\] _04023_ vssd1
+ vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__and2_1
XANTENNA__09728__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08936__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14159_ _03948_ net907 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[8\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08400__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout609 _04320_ vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08720_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[22\]
+ net842 net761 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[22\]
+ _04792_ vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_47_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_17918_ clknet_leaf_51_wb_clk_i _00002_ _01614_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.wishbone.curr_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08279__A net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1180 net1181 vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09361__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1191 net1194 vssd1 vssd1 vccd1 vccd1 net1191 sky130_fd_sc_hd__buf_4
X_08651_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[23\]
+ net642 net613 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[23\]
+ _04720_ vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__a221o_1
X_17849_ clknet_leaf_103_wb_clk_i _03192_ _01545_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[95\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_157_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08582_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[25\]
+ net753 net734 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09113__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08467__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13124__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11433__A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09203_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[10\]
+ net715 _05252_ _05255_ vssd1 vssd1 vccd1 vccd1 _05256_ sky130_fd_sc_hd__o22a_4
XFILLER_0_57_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12963__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout325_A net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14744__A net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10049__A net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09134_ _05186_ _05187_ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__or2_2
XFILLER_0_44_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12420__A0 _03612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09065_ _04158_ _04353_ _04157_ vssd1 vssd1 vccd1 vccd1 _05124_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1234_A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14182__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold630 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2044 sky130_fd_sc_hd__dlygate4sd3_1
Xhold641 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2055 sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[63\] vssd1 vssd1
+ vccd1 vccd1 net2066 sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2077 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold674 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2088 sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[15\] vssd1 vssd1
+ vccd1 vccd1 net2099 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1022_X net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_196_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold696 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[2\] vssd1
+ vssd1 vccd1 vccd1 net2110 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09967_ _05927_ _05995_ vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout861_A _04296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout482_X net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08918_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[16\]
+ net617 net598 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[16\]
+ _04982_ vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__a221o_1
X_09898_ _04513_ _04514_ vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__nor2_2
Xhold1330 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2744 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09723__D net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1341 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net2755 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1352 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2766 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_86_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08849_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[18\]
+ net782 _04916_ net853 vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__a211o_1
Xhold1363 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2777 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1374 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 net2788 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout747_X net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1385 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net2799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1396 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net2810 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11860_ _07669_ _07671_ vssd1 vssd1 vccd1 vccd1 _07672_ sky130_fd_sc_hd__and2_1
XANTENNA__09104__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10811_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[15\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06808_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11791_ _07587_ _07589_ vssd1 vssd1 vccd1 vccd1 _07603_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout914_X net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12439__A _07840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08458__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13034__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13530_ net2741 net221 net403 vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10742_ _05735_ net511 net334 _06298_ _06740_ vssd1 vssd1 vccd1 vccd1 _06741_ sky130_fd_sc_hd__o221a_1
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10673_ _04158_ _05506_ vssd1 vssd1 vccd1 vccd1 _06676_ sky130_fd_sc_hd__nor2_1
X_13461_ net200 net2079 net410 vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__mux2_1
XANTENNA__12873__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_173_Right_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15200_ net1103 vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__inv_2
X_12412_ _03657_ net1897 net214 vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__mux2_1
X_16180_ net1153 vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13392_ net2684 net325 net423 vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__mux2_1
XANTENNA__11489__S net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15131_ net1176 vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__inv_2
X_12343_ _08022_ _03518_ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10973__A0 _06464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08630__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12274_ _03564_ _03566_ vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__and2_1
X_15062_ net1084 vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_79_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08918__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11225_ net1670 net731 _07188_ vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__o21a_1
X_14013_ team_05_WB.instance_to_wrap.CPU_DAT_O\[6\] net546 _07451_ vssd1 vssd1 vccd1
+ vccd1 _03883_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11156_ _07075_ _07093_ vssd1 vssd1 vccd1 vccd1 _07122_ sky130_fd_sc_hd__nand2_2
XANTENNA__13717__B _06464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13209__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10107_ _06133_ _06134_ vssd1 vssd1 vccd1 vccd1 _06135_ sky130_fd_sc_hd__nand2_1
X_11087_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[1\] _04164_
+ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[2\] vssd1 vssd1
+ vccd1 vccd1 _07054_ sky130_fd_sc_hd__a21oi_1
X_15964_ net1299 vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__inv_2
X_17703_ clknet_leaf_86_wb_clk_i _03046_ _01399_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[77\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09343__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09770__X _05801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14915_ net1205 vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10038_ _04491_ _05770_ vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__nor2_1
X_15895_ net1292 vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_125_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13733__A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17634_ clknet_leaf_70_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[1\]
+ _01330_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14846_ net1066 vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17565_ clknet_leaf_113_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[2\]
+ _01261_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_14777_ net1051 vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__inv_2
XANTENNA__08449__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11989_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[21\] net995 net356
+ _07800_ net548 vssd1 vssd1 vccd1 vccd1 _07801_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_59_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16516_ clknet_leaf_183_wb_clk_i _02146_ _00212_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_173_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13728_ net905 _06219_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[28\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_14_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_173_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17496_ clknet_leaf_42_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[31\]
+ _01192_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_165_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_165_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_129_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16447_ clknet_leaf_155_wb_clk_i _02077_ _00143_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12783__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13659_ net2045 net197 net385 vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_140_Right_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16378_ clknet_leaf_30_wb_clk_i _02008_ _00074_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18117_ clknet_leaf_46_wb_clk_i _00031_ _01813_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15329_ net1224 vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18048_ net1037 _03386_ _01744_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_1_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08909__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10716__B1 _04275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout406 net407 vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__clkbuf_8
X_09821_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[20\]
+ net648 net640 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[20\]
+ _05851_ vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__a221o_1
Xfanout417 _03726_ vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__clkbuf_4
Xfanout428 net431 vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__buf_6
Xfanout439 _03721_ vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__buf_4
XANTENNA__13119__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09752_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[0\]
+ net886 net868 net861 vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_33_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09334__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08703_ _04772_ _04773_ _04774_ _04775_ vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__or4_1
XANTENNA__14326__A1_N net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12958__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09683_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[1\]
+ net878 net872 net864 vssd1 vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__and4_1
XANTENNA__08688__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08634_ _04702_ _04706_ _04707_ _04708_ vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__or4_1
X_08565_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[25\]
+ net669 net596 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[25\]
+ _04640_ vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_81_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout442_A _03716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1184_A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14177__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12641__A0 _03650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08496_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[27\]
+ net827 net746 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12693__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14474__A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08860__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout707_A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09117_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[12\]
+ net850 net841 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[12\]
+ _05172_ vssd1 vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08612__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09718__D _04418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09048_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[13\]
+ net682 net610 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout697_X net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold460 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[74\] vssd1 vssd1
+ vccd1 vccd1 net1874 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10707__A0 _06706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold471 _00004_ vssd1 vssd1 vccd1 vccd1 net1885 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12612__D_N _03659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11010_ net963 _06591_ _06985_ vssd1 vssd1 vccd1 vccd1 _06986_ sky130_fd_sc_hd__a21oi_1
Xhold482 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[23\] vssd1 vssd1
+ vccd1 vccd1 net1896 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold493 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[108\] vssd1 vssd1
+ vccd1 vccd1 net1907 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout864_X net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout940 net943 vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__buf_2
XANTENNA__13029__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout951 _04363_ vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__clkbuf_2
Xfanout962 net964 vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__buf_2
Xfanout973 net977 vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout984 _03763_ vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__clkbuf_2
Xfanout995 _07470_ vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12961_ net306 net2498 net468 vssd1 vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__mux2_1
XANTENNA__08679__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12868__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1160 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1171 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net2585 sky130_fd_sc_hd__dlygate4sd3_1
X_14700_ net1077 vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__inv_2
X_11912_ _07529_ _07723_ vssd1 vssd1 vccd1 vccd1 _07724_ sky130_fd_sc_hd__nor2_1
Xhold1182 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net2596 sky130_fd_sc_hd__dlygate4sd3_1
X_15680_ net1150 vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_142_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12880__A0 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1193 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net2607 sky130_fd_sc_hd__dlygate4sd3_1
X_12892_ net325 net2094 net476 vssd1 vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ net1105 vssd1 vssd1 vccd1 vccd1 _00261_ sky130_fd_sc_hd__inv_2
X_11843_ _07653_ _07654_ vssd1 vssd1 vccd1 vccd1 _07655_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09628__B2 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12632__A0 _03664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17350_ clknet_leaf_34_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[14\]
+ _01046_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14562_ net1217 vssd1 vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11774_ _07565_ _07569_ _07571_ vssd1 vssd1 vccd1 vccd1 _07586_ sky130_fd_sc_hd__and3_1
X_16301_ net1154 vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13513_ net2108 net280 net404 vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__mux2_1
X_17281_ clknet_leaf_149_wb_clk_i _02911_ _00977_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10725_ net512 _06723_ _06724_ vssd1 vssd1 vccd1 vccd1 _06725_ sky130_fd_sc_hd__o21a_1
X_14493_ net1092 vssd1 vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08851__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16232_ net1215 vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__inv_2
X_13444_ net2262 net272 net412 vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10656_ _06379_ net347 vssd1 vssd1 vccd1 vccd1 _06660_ sky130_fd_sc_hd__or2_1
XANTENNA__11199__B1 _07120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17468__Q team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16163_ net1163 vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__inv_2
Xclkload16 clknet_leaf_201_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload16/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_3_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13375_ net2152 net266 net420 vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__mux2_1
Xclkload27 clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload27/Y sky130_fd_sc_hd__inv_6
X_10587_ net513 _06134_ _06136_ _06594_ vssd1 vssd1 vccd1 vccd1 _06595_ sky130_fd_sc_hd__a31o_1
XFILLER_0_23_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload38 clknet_leaf_187_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload38/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_118_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload49 clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload49/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_140_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15114_ net1111 vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__inv_2
X_12326_ _03531_ _03536_ _03540_ net355 _07924_ vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__a32o_1
X_16094_ net1309 vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10136__B net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13728__A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09159__A3 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15045_ net1196 vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__inv_2
X_12257_ _03512_ _03543_ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__nor2_1
XANTENNA__09013__C1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16104__A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11208_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[117\] _07103_
+ _07106_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[21\] vssd1 vssd1
+ vccd1 vccd1 _07172_ sky130_fd_sc_hd__a22o_1
XANTENNA__14125__A2_N net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12188_ _07987_ _07995_ _07998_ vssd1 vssd1 vccd1 vccd1 _08000_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_166_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09644__C net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11139_ _07076_ _07087_ vssd1 vssd1 vccd1 vccd1 _07105_ sky130_fd_sc_hd__nor2_4
X_16996_ clknet_leaf_194_wb_clk_i _02626_ _00692_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09316__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15947_ net1304 vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__inv_2
XANTENNA__12778__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17580__D team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[17\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15878_ net1267 vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__inv_2
XANTENNA__08557__A _04613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17617_ clknet_leaf_49_wb_clk_i _02988_ _01313_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_14829_ net1081 vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08350_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[30\]
+ net638 net622 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__a22o_1
X_17548_ clknet_leaf_50_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[19\]
+ _01244_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12623__A0 _03610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09095__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08281_ _04236_ _04240_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[24\]
+ _04230_ vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__o211a_1
X_17479_ clknet_leaf_37_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[14\]
+ _01175_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08842__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13402__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14376__B1 _07451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11430__B team_05_WB.instance_to_wrap.wishbone.curr_state\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_62_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_112_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout203 net204 vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__buf_4
Xfanout214 net215 vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__buf_4
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout225 _06271_ vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout392_A _03732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout236 net237 vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__clkbuf_2
X_09804_ _05104_ _05834_ _05102_ vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__a21o_1
Xfanout247 net249 vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__buf_2
Xfanout258 _06442_ vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_31_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout269 _06499_ vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_66_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09735_ net587 _05757_ _05758_ net586 vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__and4_1
XFILLER_0_158_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10997__A _04170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout657_A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09570__B net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09666_ net571 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[1\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[1\] vssd1 vssd1 vccd1
+ vccd1 _05699_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13804__C net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08617_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[24\]
+ net669 net626 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout445_X net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09597_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[2\]
+ net591 _05628_ _05632_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[2\]
+ sky130_fd_sc_hd__o22a_4
XANTENNA_fanout824_A net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1187_X net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12614__A0 _03661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08548_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[26\]
+ net800 net762 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__a22o_1
XANTENNA__09086__A2 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08294__B1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[21\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout612_X net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08479_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[27\]
+ net634 net612 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08473__Y _04552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13312__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10510_ net888 _06521_ _06520_ net554 vssd1 vssd1 vccd1 vccd1 _06522_ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11490_ _07346_ _07400_ vssd1 vssd1 vccd1 vccd1 _07401_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10441_ _06446_ _06456_ _04275_ vssd1 vssd1 vccd1 vccd1 _06457_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_98_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18404__A net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10372_ net1020 _05885_ net552 vssd1 vssd1 vccd1 vccd1 _06391_ sky130_fd_sc_hd__a21oi_1
X_13160_ _04253_ _04257_ net562 vssd1 vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__or3_4
XANTENNA_fanout981_X net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12111_ net547 _07622_ vssd1 vssd1 vccd1 vccd1 _07923_ sky130_fd_sc_hd__nand2_2
Xclkbuf_4_10__f_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_10__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_13091_ net323 net2850 net453 vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12042_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[27\] team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[29\]
+ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[30\] net993 vssd1 vssd1
+ vccd1 vccd1 _07854_ sky130_fd_sc_hd__o31a_1
XANTENNA__09546__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold290 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[111\] vssd1 vssd1
+ vccd1 vccd1 net1704 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_72_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09010__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16850_ clknet_leaf_135_wb_clk_i _02480_ _00546_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_144_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15801_ net1276 vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__inv_2
Xfanout770 _04407_ vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__clkbuf_8
Xfanout781 _04403_ vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__buf_4
X_16781_ clknet_leaf_160_wb_clk_i _02411_ _00477_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout792 net793 vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__buf_4
XANTENNA__12598__S net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13993_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[11\] net980 vssd1
+ vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15732_ net1305 vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12944_ net260 net2610 net471 vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15663_ net1158 vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__inv_2
X_12875_ net263 net2756 net476 vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__mux2_1
X_17402_ clknet_leaf_69_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[2\]
+ _01098_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_14614_ net1091 vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__inv_2
X_18382_ net1367 vssd1 vssd1 vccd1 vccd1 la_data_out[30] sky130_fd_sc_hd__buf_2
X_11826_ _07637_ vssd1 vssd1 vccd1 vccd1 _07638_ sky130_fd_sc_hd__inv_2
XANTENNA__09077__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15594_ net1283 vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__inv_2
X_17333_ clknet_leaf_71_wb_clk_i _02963_ _01029_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13730__B _06108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14545_ net1189 vssd1 vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__inv_2
X_11757_ _07565_ _07566_ _07563_ _07564_ vssd1 vssd1 vccd1 vccd1 _07569_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_166_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08824__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10631__A2 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17264_ clknet_leaf_151_wb_clk_i _02894_ _00960_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10708_ net554 _06708_ vssd1 vssd1 vccd1 vccd1 _06709_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14476_ net1111 vssd1 vssd1 vccd1 vccd1 _00106_ sky130_fd_sc_hd__inv_2
X_11688_ net59 net60 vssd1 vssd1 vccd1 vccd1 _07502_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09639__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16215_ net1243 vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload105 clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload105/Y sky130_fd_sc_hd__bufinv_16
X_13427_ _04252_ net557 _03701_ vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__and3_4
X_10639_ net1021 _05421_ net552 _06643_ vssd1 vssd1 vccd1 vccd1 _06644_ sky130_fd_sc_hd__o31a_1
X_17195_ clknet_leaf_188_wb_clk_i _02825_ _00891_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload116 clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload116/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_107_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload127 clknet_leaf_173_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload127/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload138 clknet_leaf_148_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload138/X sky130_fd_sc_hd__clkbuf_8
X_16146_ net1263 vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__inv_2
Xclkload149 clknet_leaf_134_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload149/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_122_840 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13358_ net321 net2842 net424 vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_168_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17575__D team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[12\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12309_ net544 _07536_ _08022_ _03516_ _03603_ vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__o32a_2
XFILLER_0_11_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16077_ net1262 vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13289_ net315 net2898 net435 vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__mux2_1
XANTENNA_wire360_A _05860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15028_ net1073 vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09001__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15673__A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput3 DAT_I[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
X_16979_ clknet_leaf_170_wb_clk_i _02609_ _00675_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_09520_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[3\]
+ net826 net745 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_180_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_180_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_18405__1374 vssd1 vssd1 vccd1 vccd1 _18405__1374/HI net1374 sky130_fd_sc_hd__conb_1
XFILLER_0_79_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09451_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[5\]
+ net831 net824 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[5\]
+ _05492_ vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08402_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[29\]
+ net686 net648 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__a22o_1
X_09382_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[6\]
+ net677 net626 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05427_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09068__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08333_ net950 net931 net929 vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__and3_1
XANTENNA__08815__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13132__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11441__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08264_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[23\] team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__nor2_2
XFILLER_0_34_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08195_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[29\] team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[28\]
+ _04277_ vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__nor3_1
XANTENNA__09225__C1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12971__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout405_A net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09240__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_93_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11159__Y _07125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1009 net1010 vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__buf_2
XANTENNA_fanout774_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout395_X net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09852__Y _05881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13307__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11616__A team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[12\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09718_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[0\]
+ net945 net938 _04418_ vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__and4_1
X_10990_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[14\] net566 _06968_
+ _06969_ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09649_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[1\]
+ net1016 net942 net932 vssd1 vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout827_X net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14927__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[29\]
+ net342 vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09059__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08925__A _04989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11611_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[15\] net995 vssd1
+ vssd1 vccd1 vccd1 _07476_ sky130_fd_sc_hd__and2_2
XFILLER_0_93_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12591_ _03620_ net1805 net203 vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__mux2_1
XANTENNA__08806__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13042__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14330_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[2\] net523
+ vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11542_ _07353_ _07444_ vssd1 vssd1 vccd1 vccd1 _07453_ sky130_fd_sc_hd__nor2_1
XFILLER_0_167_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10238__Y _06263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14261_ _04020_ _04044_ vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11473_ _07353_ _07383_ vssd1 vssd1 vccd1 vccd1 _07384_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12881__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14662__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16000_ net1112 vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__inv_2
XANTENNA_input70_A wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13212_ _06554_ net2821 net350 vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__mux2_1
X_10424_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[19\] net904 net968
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[19\] _06440_ vssd1
+ vssd1 vccd1 vccd1 _06441_ sky130_fd_sc_hd__a221o_1
XFILLER_0_122_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14192_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[4\] _03998_
+ vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11497__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13143_ net267 net2911 net444 vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__mux2_1
X_10355_ net337 _06140_ _06156_ net333 _06374_ vssd1 vssd1 vccd1 vccd1 _06375_ sky130_fd_sc_hd__o221a_1
XFILLER_0_103_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09519__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17951_ clknet_leaf_43_wb_clk_i _03290_ _01647_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13074_ net257 net2666 net452 vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__mux2_1
X_10286_ _06200_ _06209_ net524 vssd1 vssd1 vccd1 vccd1 _06309_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_163_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15493__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12025_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[19\] net996 _07747_
+ net548 vssd1 vssd1 vccd1 vccd1 _07837_ sky130_fd_sc_hd__a211o_1
X_16902_ clknet_leaf_115_wb_clk_i _02532_ _00598_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_17882_ clknet_leaf_98_wb_clk_i _03225_ _01578_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13725__B _06918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16833_ clknet_leaf_148_wb_clk_i _02463_ _00529_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12330__D_N _03610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16764_ clknet_leaf_158_wb_clk_i _02394_ _00460_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13976_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[13\] _03847_ vssd1
+ vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11629__B2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09641__D net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09298__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_24_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15715_ net1142 vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__inv_2
X_12927_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[9\] _04254_
+ vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__nor2_1
XANTENNA__10301__A1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16695_ clknet_leaf_145_wb_clk_i _02325_ _00391_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15646_ net1248 vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__inv_2
X_12858_ net321 net2361 net483 vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18365_ net1350 vssd1 vssd1 vccd1 vccd1 la_data_out[13] sky130_fd_sc_hd__buf_2
X_11809_ _07606_ _07609_ _07620_ _07604_ vssd1 vssd1 vccd1 vccd1 _07621_ sky130_fd_sc_hd__o22ai_4
X_15577_ net1246 vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__inv_2
X_12789_ net309 net2816 net488 vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_1_Left_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17316_ clknet_leaf_184_wb_clk_i _02946_ _01012_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_14528_ net1195 vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18296_ net1388 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
XFILLER_0_160_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17247_ clknet_leaf_152_wb_clk_i _02877_ _00943_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12791__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14459_ net1098 vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17178_ clknet_leaf_11_wb_clk_i _02808_ _00874_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09222__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14291__B team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[27\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16129_ net1277 vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08951_ _05012_ _05013_ vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__nor2_1
XANTENNA__11317__B1 _07108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_63_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08882_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[17\]
+ net846 net795 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09289__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09503_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[4\]
+ net688 net599 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08497__B1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12966__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09694__C1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1097_A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09434_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[5\]
+ net658 net650 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12045__A1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[31\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08249__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09365_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[7\]
+ net761 net754 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[7\]
+ _05410_ vssd1 vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__a221o_1
XANTENNA__10486__S net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1264_A net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11253__C1 _07031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08316_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[31\]
+ net803 net799 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[31\]
+ _04397_ vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_502 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09296_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[8\]
+ net696 net670 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[8\]
+ _05344_ vssd1 vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__a221o_1
XANTENNA__09461__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08247_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[31\]
+ net713 net673 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[31\]
+ _04329_ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_95_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout408_X net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08178_ _04250_ _04251_ vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout891_A _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09213__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11020__A2 _06623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18287__1379 vssd1 vssd1 vccd1 vccd1 net1379 _18287__1379/LO sky130_fd_sc_hd__conb_1
X_10140_ net378 net363 vssd1 vssd1 vccd1 vccd1 _06168_ sky130_fd_sc_hd__nand2_1
Xoutput170 net170 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__clkbuf_4
XANTENNA__11308__B1 _07126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput181 net181 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout777_X net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10071_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[25\] team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[24\]
+ _06099_ vssd1 vssd1 vccd1 vccd1 _06100_ sky130_fd_sc_hd__and3_1
XANTENNA__09742__C _04287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout944_X net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13037__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13830_ net1466 net582 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[8\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_98_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13761_ net921 _06185_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[29\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08488__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10973_ _06464_ _06955_ net956 vssd1 vssd1 vccd1 vccd1 _06956_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12876__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15500_ net1164 vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_67_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12712_ net279 net2404 net496 vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__mux2_1
X_16480_ clknet_leaf_132_wb_clk_i _02110_ _00176_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13692_ net1049 _06772_ _07350_ vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_139_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_108_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15431_ net1123 vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__inv_2
X_12643_ _03641_ net1825 net202 vssd1 vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10249__X _06273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09437__C1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18150_ clknet_leaf_200_wb_clk_i _03453_ _01846_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_156_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15362_ net1226 vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11512__C _07422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12574_ net1628 _07836_ _03678_ vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_156_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09452__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17101_ clknet_leaf_159_wb_clk_i _02731_ _00797_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14313_ _04944_ _04965_ vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__and2_1
X_18081_ clknet_leaf_83_wb_clk_i _00008_ _01777_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11525_ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[26\] _07435_ net1001
+ vssd1 vssd1 vccd1 vccd1 _07436_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15293_ net1089 vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__inv_2
XANTENNA__08660__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13500__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17032_ clknet_leaf_1_wb_clk_i _02662_ _00728_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14244_ _04026_ _04032_ vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__nor2_1
X_11456_ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[2\] _07366_ net1002
+ vssd1 vssd1 vccd1 vccd1 _07367_ sky130_fd_sc_hd__mux2_2
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10407_ _05840_ _05931_ vssd1 vssd1 vccd1 vccd1 _06424_ sky130_fd_sc_hd__xnor2_4
X_14175_ net1974 net506 net909 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[24\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__08412__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11387_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[13\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[12\]
+ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[11\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[10\]
+ vssd1 vssd1 vccd1 vccd1 _07318_ sky130_fd_sc_hd__or4_1
XFILLER_0_22_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13126_ net305 net2002 net449 vssd1 vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__mux2_1
X_10338_ _06260_ _06358_ net531 vssd1 vssd1 vccd1 vccd1 _06359_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_119_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_119_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_17934_ clknet_leaf_34_wb_clk_i _03273_ _01630_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13057_ net310 net2227 net457 vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__mux2_1
X_10269_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[26\] net904 net968
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[26\] _06292_ vssd1
+ vssd1 vccd1 vccd1 _06293_ sky130_fd_sc_hd__a221o_1
X_12008_ _07765_ _07767_ _07769_ _07773_ vssd1 vssd1 vccd1 vccd1 _07820_ sky130_fd_sc_hd__or4_1
XFILLER_0_79_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17865_ clknet_leaf_100_wb_clk_i _03208_ _01561_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09652__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_147_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16816_ clknet_leaf_123_wb_clk_i _02446_ _00512_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_128_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17796_ clknet_leaf_77_wb_clk_i _03139_ _01492_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13959_ _04160_ _03830_ vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__and2_1
X_16747_ clknet_leaf_186_wb_clk_i _02377_ _00443_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08479__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12786__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16678_ clknet_leaf_115_wb_clk_i _02308_ _00374_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09691__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15629_ net1245 vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11235__C1 _07031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09948__X _05977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09150_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[11\]
+ net707 net683 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[11\]
+ _05192_ vssd1 vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__a221o_1
XFILLER_0_84_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18348_ net37 vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08101_ net1030 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__and2b_1
XFILLER_0_72_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15398__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18279_ clknet_leaf_50_wb_clk_i net1885 _01973_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instr_fetch
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11250__A2 _07119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08651__B1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09081_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[13\]
+ net778 _05138_ net854 vssd1 vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__a211o_1
XFILLER_0_114_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13410__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08032_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[17\] vssd1
+ vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__inv_2
Xinput50 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_1
Xinput61 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_1
Xinput72 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__clkbuf_1
Xhold801 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 net2215 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold812 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2226 sky130_fd_sc_hd__dlygate4sd3_1
Xhold823 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 net2237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold834 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2248 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08403__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold845 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2259 sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 net2270 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_186_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold867 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2281 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold878 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold889 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net2303 sky130_fd_sc_hd__dlygate4sd3_1
X_09983_ _06010_ _06011_ vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08934_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[16\]
+ net829 net760 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1501 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 net2915 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1512 team_05_WB.instance_to_wrap.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 net2926
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08865_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[17\]
+ net695 net651 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout472_A _03706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1523 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 net2937 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1534 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2948 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1545 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 net2959 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1556 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[6\] vssd1
+ vssd1 vccd1 vccd1 net2970 sky130_fd_sc_hd__dlygate4sd3_1
X_08796_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[19\]
+ net833 net764 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[19\]
+ _04863_ vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_88_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12696__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_154_Right_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08746__Y _04818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout737_A net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_64_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13812__C net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12018__A1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[20\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09417_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[6\]
+ net779 _05458_ _05460_ net855 vssd1 vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13215__A0 _06605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout904_A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08890__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08194__B team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[26\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09348_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[7\]
+ net649 net634 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[7\]
+ _05384_ vssd1 vssd1 vccd1 vccd1 _05395_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09434__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11241__A2 _07106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09279_ _05315_ _05324_ _05328_ net592 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[9\]
+ sky130_fd_sc_hd__o32a_4
XFILLER_0_90_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12725__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13320__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11310_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[40\] _07113_
+ _07118_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[64\] vssd1 vssd1
+ vccd1 vccd1 _07269_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_151_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12290_ _03580_ _03582_ _03584_ _03577_ vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_151_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout894_X net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11241_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[20\] _07106_
+ _07109_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[76\] _07190_
+ vssd1 vssd1 vccd1 vccd1 _07204_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_73_Left_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11172_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[63\] _07115_
+ _07121_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[87\] _07137_
+ vssd1 vssd1 vccd1 vccd1 _07138_ sky130_fd_sc_hd__a221o_1
XFILLER_0_140_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10123_ _06149_ _06150_ vssd1 vssd1 vccd1 vccd1 _06151_ sky130_fd_sc_hd__nand2_1
X_15980_ net1169 vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input33_A DAT_I[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10054_ _06003_ _06033_ _06082_ vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__o21ai_1
X_14931_ net1212 vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__inv_2
X_17650_ clknet_leaf_54_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[17\]
+ _01346_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14862_ net1179 vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__inv_2
X_13813_ net1568 net974 net723 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[24\]
+ sky130_fd_sc_hd__and3_1
X_16601_ clknet_leaf_9_wb_clk_i _02231_ _00297_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17581_ clknet_leaf_72_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[18\]
+ _01277_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_82_Left_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14793_ net1215 vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_158_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16532_ clknet_leaf_120_wb_clk_i _02162_ _00228_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_158_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13744_ net922 _06557_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[12\]
+ sky130_fd_sc_hd__nor2_1
X_10956_ net1042 _06940_ _06941_ net961 vssd1 vssd1 vccd1 vccd1 _06942_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_123_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16463_ clknet_leaf_134_wb_clk_i _02093_ _00159_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13675_ net2367 net271 net384 vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__mux2_1
XANTENNA__08881__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10887_ _06779_ _06883_ vssd1 vssd1 vccd1 vccd1 _06884_ sky130_fd_sc_hd__and2_1
XFILLER_0_167_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15414_ net1138 vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__inv_2
X_18202_ clknet_leaf_37_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[23\]
+ _01897_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12626_ _03614_ net1759 net202 vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16394_ clknet_leaf_3_wb_clk_i _02024_ _00090_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09425__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10139__B net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18133_ clknet_leaf_47_wb_clk_i _00029_ _01829_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_15345_ net1188 vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__inv_2
X_12557_ _03620_ net1787 net207 vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__mux2_1
XANTENNA__11232__A2 _07091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08633__B1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13230__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11508_ _07414_ _07418_ _07416_ _07412_ vssd1 vssd1 vccd1 vccd1 _07419_ sky130_fd_sc_hd__or4bb_1
X_18064_ clknet_leaf_98_wb_clk_i _03402_ _01760_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_91_Left_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15276_ net1077 vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12488_ net1655 _03620_ _03674_ vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__mux2_1
XANTENNA__09647__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold108 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[29\] vssd1 vssd1
+ vccd1 vccd1 net1522 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17015_ clknet_leaf_144_wb_clk_i _02645_ _00711_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_14227_ team_05_WB.instance_to_wrap.total_design.keypad0.counter\[10\] team_05_WB.instance_to_wrap.total_design.keypad0.counter\[11\]
+ _04022_ vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__and3_1
Xhold119 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[9\]
+ vssd1 vssd1 vccd1 vccd1 net1533 sky130_fd_sc_hd__dlygate4sd3_1
X_11439_ _07349_ _07351_ team_05_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 _07352_ sky130_fd_sc_hd__o21a_2
XFILLER_0_106_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14158_ _03930_ net907 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[7\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17583__D team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[20\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13109_ net259 net2344 net449 vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__mux2_1
X_14089_ _03954_ _03955_ vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17917_ clknet_leaf_51_wb_clk_i _00001_ _01613_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.wishbone.curr_state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11299__A2 _07116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12496__A1 _03604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08279__B team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[21\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1170 net1175 vssd1 vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__buf_2
Xfanout1181 net1186 vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__buf_2
X_08650_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[23\]
+ net709 net639 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[23\]
+ _04723_ vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__a221o_1
X_17848_ clknet_leaf_90_wb_clk_i _03191_ _01544_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[94\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1192 net1194 vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__buf_4
XFILLER_0_89_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08581_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[25\]
+ net819 net775 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_87_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_17779_ clknet_leaf_89_wb_clk_i _03122_ _01475_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14297__A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13405__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_16_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11433__B net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18286__1378 vssd1 vssd1 vccd1 vccd1 net1378 _18286__1378/LO sky130_fd_sc_hd__conb_1
XFILLER_0_14_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09202_ _05239_ _05242_ _05244_ _05254_ vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__or4_1
XFILLER_0_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09416__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09133_ _05187_ vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11223__A2 _07116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09397__Y _05442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08624__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout220_A net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13140__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout318_A _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09064_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[13\]
+ net716 _05116_ _05122_ vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_103_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold620 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net2034 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold631 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2045 sky130_fd_sc_hd__dlygate4sd3_1
Xhold642 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2056 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1227_A net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold653 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2067 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09854__A _05881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold664 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2078 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10195__C1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold675 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net2089 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold686 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 net2100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2111 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout687_A net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09966_ _05909_ _05993_ _05916_ vssd1 vssd1 vccd1 vccd1 _05995_ sky130_fd_sc_hd__a21boi_1
XANTENNA__09573__B net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13807__C net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1015_X net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08917_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[16\]
+ net668 net614 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__a22o_1
XANTENNA__12487__A1 _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09897_ net380 _04466_ vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_85_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1320 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2734 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout854_A _04367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout475_X net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09352__A1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[19\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1331 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net2745 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09352__B2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[27\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10004__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08848_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[18\]
+ net802 net748 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__a22o_1
Xhold1342 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2756 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1353 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1364 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net2778 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1375 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2789 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1386 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2800 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13823__B net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08779_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[19\]
+ net687 net601 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout642_X net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1397 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2811 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13315__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10810_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[16\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06807_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_0_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ net549 _07600_ vssd1 vssd1 vccd1 vccd1 _07602_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09655__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10741_ _05734_ _06739_ vssd1 vssd1 vccd1 vccd1 _06740_ sky130_fd_sc_hd__nand2_1
XANTENNA__08863__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13460_ team_05_WB.instance_to_wrap.total_design.core.instr_fetch _04258_ _04261_
+ _03708_ vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__or4_4
X_10672_ net890 _06672_ _06674_ net555 vssd1 vssd1 vccd1 vccd1 _06675_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_153_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09407__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12411_ net1772 _07791_ _03667_ vssd1 vssd1 vccd1 vccd1 _03219_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11214__A2 _07101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12411__A1 _07791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08615__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13391_ net1925 net323 net423 vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__mux2_1
XANTENNA__13050__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15130_ net1055 vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12342_ _07658_ _03616_ _03636_ _03541_ vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__o22a_1
XFILLER_0_106_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15061_ net1059 vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__inv_2
X_12273_ _03563_ _03567_ _03564_ vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__o21ai_1
XANTENNA__14670__A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14012_ _03798_ _03882_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[5\]
+ sky130_fd_sc_hd__nor2_1
X_11224_ _07177_ _07179_ _07182_ _07187_ vssd1 vssd1 vccd1 vccd1 _07188_ sky130_fd_sc_hd__or4_1
XANTENNA__08394__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11155_ _07094_ _07114_ vssd1 vssd1 vccd1 vccd1 _07121_ sky130_fd_sc_hd__nor2_4
XFILLER_0_105_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10106_ _05123_ net361 vssd1 vssd1 vccd1 vccd1 _06134_ sky130_fd_sc_hd__nand2_1
XANTENNA__12478__A1 _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11086_ _07032_ _07034_ _07044_ _07040_ vssd1 vssd1 vccd1 vccd1 _07053_ sky130_fd_sc_hd__a31oi_1
X_15963_ net1304 vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__inv_2
XANTENNA__10489__A0 _06500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17702_ clknet_leaf_87_wb_clk_i _03045_ _01398_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[76\]
+ sky130_fd_sc_hd__dfrtp_1
X_14914_ net1228 vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__inv_2
X_10037_ _04428_ net510 _06060_ net336 _06053_ vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__o221a_1
X_15894_ net1256 vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_125_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_125_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13733__B _06743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17633_ clknet_leaf_70_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[0\]
+ _01329_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14845_ net1089 vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__inv_2
XFILLER_0_172_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15006__A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14776_ net1242 vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__inv_2
X_17564_ clknet_leaf_114_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[1\]
+ _01260_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11988_ _07777_ _07785_ _07795_ vssd1 vssd1 vccd1 vccd1 _07800_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13727_ net900 _06907_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[27\]
+ sky130_fd_sc_hd__nor2_1
X_16515_ clknet_leaf_198_wb_clk_i _02145_ _00211_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10939_ _06791_ _06792_ vssd1 vssd1 vccd1 vccd1 _06928_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_173_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17495_ clknet_leaf_36_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[30\]
+ _01191_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16446_ clknet_leaf_185_wb_clk_i _02076_ _00142_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13658_ _04256_ _04259_ _03697_ vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17578__D team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[15\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11540__Y _07451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12609_ _03641_ net1853 net204 vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12402__A1 _03641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08606__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16377_ clknet_leaf_9_wb_clk_i _02007_ _00073_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13589_ net2462 net322 net397 vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18116_ clknet_leaf_46_wb_clk_i _00021_ _01812_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_15328_ net1102 vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10156__Y _06184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_134_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_134_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18047_ net1038 _03385_ _01743_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_15259_ net1176 vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__inv_2
XANTENNA__08385__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09820_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[20\]
+ net668 net652 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__a22o_1
Xfanout407 _03729_ vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__buf_4
Xfanout418 net419 vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11709__A _07476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout429 net431 vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_129_Left_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09751_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[0\]
+ net887 net863 net859 vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__and4_1
XANTENNA__12469__A1 _03650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08702_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[22\]
+ net667 net650 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[22\]
+ _04759_ vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__a221o_1
XFILLER_0_146_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09682_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[1\]
+ net883 net874 net862 vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__and4_1
X_08633_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[24\]
+ net843 net827 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[24\]
+ _04700_ vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout268_A _06499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13135__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09098__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08564_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[25\]
+ net657 net634 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_81_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08845__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12974__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08495_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[27\]
+ net717 _04568_ _04572_ vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__o22ai_4
XANTENNA_fanout435_A _03722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1177_A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_138_Left_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout602_A net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09568__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09116_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[12\]
+ net829 net745 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09270__B1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09047_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[13\]
+ net703 net655 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold450 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[115\] vssd1 vssd1
+ vccd1 vccd1 net1864 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09022__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold461 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[53\] vssd1 vssd1
+ vccd1 vccd1 net1875 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout592_X net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold472 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[47\] vssd1 vssd1
+ vccd1 vccd1 net1886 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_147_Left_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08376__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold483 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[57\] vssd1 vssd1
+ vccd1 vccd1 net1897 sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 net84 vssd1 vssd1 vccd1 vccd1 net1908 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout930 net931 vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__buf_2
Xfanout941 net943 vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__buf_1
X_09949_ _05880_ _05886_ vssd1 vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__nor2_2
Xfanout963 net964 vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__buf_2
XANTENNA_fanout857_X net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout974 net977 vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__buf_2
Xfanout985 net988 vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__buf_2
Xfanout996 _07470_ vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12960_ net326 net2036 net471 vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_5_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1150 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2564 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11911_ _07707_ _07713_ vssd1 vssd1 vccd1 vccd1 _07723_ sky130_fd_sc_hd__xnor2_1
Xhold1161 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2575 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1172 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2586 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1183 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net2597 sky130_fd_sc_hd__dlygate4sd3_1
X_12891_ net323 net2336 net476 vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__mux2_1
XANTENNA__09750__C net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1194 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2608 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13045__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14630_ net1231 vssd1 vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__inv_2
X_11842_ _07625_ _07627_ vssd1 vssd1 vccd1 vccd1 _07654_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_16_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09628__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_156_Left_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ net1236 vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__inv_2
XANTENNA__12884__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08836__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11773_ _07568_ _07571_ _07584_ _07566_ vssd1 vssd1 vccd1 vccd1 _07585_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__14665__A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16300_ net1154 vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__inv_2
X_13512_ net2777 net283 net407 vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17280_ clknet_leaf_129_wb_clk_i _02910_ _00976_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10724_ net512 _06696_ vssd1 vssd1 vccd1 vccd1 _06724_ sky130_fd_sc_hd__nand2_1
X_14492_ net1063 vssd1 vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__inv_2
X_16231_ net1220 vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__inv_2
X_13443_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[16\]
+ net267 net412 vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10655_ net890 _06658_ _06657_ net555 vssd1 vssd1 vccd1 vccd1 _06659_ sky130_fd_sc_hd__a211o_1
XFILLER_0_125_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16162_ net1164 vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13374_ net2650 net257 net420 vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload17 clknet_leaf_202_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload17/Y sky130_fd_sc_hd__inv_8
XFILLER_0_106_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09261__B1 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload28 clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload28/Y sky130_fd_sc_hd__bufinv_16
X_10586_ net516 _06126_ _06137_ vssd1 vssd1 vccd1 vccd1 _06594_ sky130_fd_sc_hd__and3_1
XANTENNA__10946__A1 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15113_ net1221 vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__inv_2
Xclkload39 clknet_leaf_188_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload39/X sky130_fd_sc_hd__clkbuf_4
X_12325_ _03609_ _03619_ vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__nand2_2
X_16093_ net1309 vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_165_Left_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15044_ net1205 vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__inv_2
X_12256_ _03550_ vssd1 vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__inv_2
XANTENNA__13728__B _06219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11207_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[45\] _07091_
+ _07110_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[53\] _07170_
+ vssd1 vssd1 vccd1 vccd1 _07171_ sky130_fd_sc_hd__a221o_1
XANTENNA__08367__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12187_ _07995_ _07998_ vssd1 vssd1 vccd1 vccd1 _07999_ sky130_fd_sc_hd__nand2_1
X_18285__1377 vssd1 vssd1 vccd1 vccd1 net1377 _18285__1377/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_166_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09644__D net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11138_ _07039_ _07076_ vssd1 vssd1 vccd1 vccd1 _07104_ sky130_fd_sc_hd__nor2_4
X_16995_ clknet_leaf_199_wb_clk_i _02625_ _00691_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13744__A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11069_ _04162_ _07035_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[5\]
+ vssd1 vssd1 vccd1 vccd1 _07036_ sky130_fd_sc_hd__a21oi_4
X_15946_ net1295 vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15877_ net1252 vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17616_ clknet_leaf_50_wb_clk_i _02987_ _01312_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14828_ net1071 vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__inv_2
XANTENNA__09619__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17547_ clknet_leaf_49_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[18\]
+ _01243_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14759_ net1242 vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08280_ net573 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[21\] vssd1
+ vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__or2_2
XFILLER_0_172_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17478_ clknet_leaf_41_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[13\]
+ _01174_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_144_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16429_ clknet_leaf_159_wb_clk_i _02059_ _00125_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09004__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10614__Y _06621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08358__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout204 _03681_ vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__buf_4
Xfanout215 _03668_ vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__buf_4
Xfanout226 net229 vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__clkbuf_2
X_09803_ _05829_ _05833_ _05146_ vssd1 vssd1 vccd1 vccd1 _05834_ sky130_fd_sc_hd__a21o_2
Xfanout237 _06346_ vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__clkbuf_2
Xfanout248 net249 vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12969__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout259 net262 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__buf_2
XANTENNA_fanout385_A net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09734_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[0\]
+ net829 _05765_ net854 vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_2_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_31_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_2_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09665_ _05692_ _05693_ _05698_ net591 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[1\]
+ sky130_fd_sc_hd__o32a_4
XANTENNA_fanout552_A net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10489__S net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09570__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1294_A net1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08616_ _04684_ _04686_ _04688_ _04690_ vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__or4_1
XANTENNA__08530__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09596_ _05623_ _05629_ _05630_ _05631_ vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__or4_1
XFILLER_0_167_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08547_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[26\]
+ net780 net750 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[26\]
+ _04623_ vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__a221o_1
XANTENNA__08818__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout340_X net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout817_A _04388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout438_X net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13820__C net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08478_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[27\]
+ net638 net630 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_838 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10077__X _06106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout605_X net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10440_ net348 _06451_ _06455_ vssd1 vssd1 vccd1 vccd1 _06456_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09243__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08597__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10371_ net892 _06387_ _06389_ vssd1 vssd1 vccd1 vccd1 _06390_ sky130_fd_sc_hd__o21a_1
XFILLER_0_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12110_ _07916_ _07918_ vssd1 vssd1 vccd1 vccd1 _07922_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_14_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13090_ net311 net2067 net452 vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__mux2_1
XANTENNA__09745__C net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10524__Y _06536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_148_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08349__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12041_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[19\] team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[20\]
+ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[21\] team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[24\]
+ net993 vssd1 vssd1 vccd1 vccd1 _07853_ sky130_fd_sc_hd__o41a_1
Xhold280 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[11\] vssd1 vssd1
+ vccd1 vccd1 net1694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[25\] vssd1 vssd1
+ vccd1 vccd1 net1705 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11353__B2 team_05_WB.instance_to_wrap.total_design.data_from_keypad\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12879__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout760 net763 vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__clkbuf_8
X_15800_ net1275 vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__inv_2
Xfanout771 _04406_ vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__clkbuf_8
Xfanout782 net785 vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__clkbuf_8
X_13992_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[11\] net980 vssd1
+ vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__or2_1
X_16780_ clknet_leaf_0_wb_clk_i _02410_ _00476_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout793 _04396_ vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__buf_4
XANTENNA__09849__A2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[19\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15731_ net1305 vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__inv_2
X_12943_ net265 net2070 net468 vssd1 vssd1 vccd1 vccd1 _02696_ sky130_fd_sc_hd__mux2_1
XANTENNA__08521__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15662_ net1140 vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__inv_2
X_12874_ net256 net2879 net477 vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__mux2_1
X_17401_ clknet_leaf_60_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[1\]
+ _01097_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14613_ net1058 vssd1 vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__inv_2
X_11825_ _07559_ _07596_ vssd1 vssd1 vccd1 vccd1 _07637_ sky130_fd_sc_hd__and2b_1
XANTENNA__12605__A1 _07821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08809__B1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[19\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18381_ net1366 vssd1 vssd1 vccd1 vccd1 la_data_out[29] sky130_fd_sc_hd__buf_2
X_15593_ net1248 vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__inv_2
XANTENNA__13503__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14310__A1_N team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[16\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14544_ net1092 vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__inv_2
X_17332_ clknet_leaf_111_wb_clk_i _02962_ _01028_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11756_ _07567_ vssd1 vssd1 vccd1 vccd1 _07568_ sky130_fd_sc_hd__inv_2
XANTENNA__09482__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14358__A1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10707_ _06706_ _06707_ net892 vssd1 vssd1 vccd1 vccd1 _06708_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17263_ clknet_leaf_141_wb_clk_i _02893_ _00959_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_14475_ net1068 vssd1 vssd1 vccd1 vccd1 _00105_ sky130_fd_sc_hd__inv_2
X_11687_ net56 net55 net58 net57 vssd1 vssd1 vccd1 vccd1 _07501_ sky130_fd_sc_hd__or4_1
XFILLER_0_126_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09639__D net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16214_ net1104 vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__inv_2
X_13426_ net1953 net307 net417 vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__mux2_1
XANTENNA__09776__X _05807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10638_ _05420_ _06051_ net510 _05423_ vssd1 vssd1 vccd1 vccd1 _06643_ sky130_fd_sc_hd__o2bb2a_1
X_17194_ clknet_leaf_196_wb_clk_i _02824_ _00890_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload106 clknet_leaf_158_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload106/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__10919__A1 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload117 clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload117/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_107_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload128 clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload128/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__14325__A1_N _05801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16145_ net1263 vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__inv_2
Xclkload139 clknet_leaf_149_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload139/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__08588__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13739__A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13357_ net312 net2662 net424 vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__mux2_1
X_10569_ _05208_ _05235_ _04158_ vssd1 vssd1 vccd1 vccd1 _06578_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_168_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12308_ net250 _03551_ _03602_ _08022_ vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_23_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16076_ net1259 vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13288_ net317 net2239 net433 vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__mux2_1
X_15027_ net1218 vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_53_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12239_ _03518_ _03519_ vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12789__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08760__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09671__B net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16978_ clknet_leaf_123_wb_clk_i _02608_ _00674_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14289__B _06185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput4 DAT_I[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
X_15929_ net1271 vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08512__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09450_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[5\]
+ net789 net758 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05492_ sky130_fd_sc_hd__a22o_1
X_08401_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[29\]
+ net672 net615 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[29\]
+ _04480_ vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__a221o_1
XFILLER_0_118_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09381_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[6\]
+ net712 net704 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[6\]
+ _05425_ vssd1 vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__a221o_1
XFILLER_0_52_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13413__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08332_ net943 net937 net928 vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09473__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10083__A1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11441__B net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11280__B1 _07106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08263_ net967 _04269_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__o21a_1
XFILLER_0_117_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_92_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08194_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[27\] team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[26\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[25\] vssd1 vssd1
+ vccd1 vccd1 _04277_ sky130_fd_sc_hd__or3_1
XFILLER_0_171_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10057__B team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout300_A _06621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1042_A net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09565__C net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1012 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12532__A0 _07797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12699__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_X net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08751__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10360__X _06380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09581__B net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09717_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[0\]
+ net950 net939 _04418_ vssd1 vssd1 vccd1 vccd1 _05749_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout555_X net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08197__B team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[30\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08503__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09648_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[1\]
+ net940 net935 net927 vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__and4_1
XANTENNA__10310__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13831__B net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout722_X net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09579_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[2\]
+ net946 net935 net932 vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__and4_1
XFILLER_0_171_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12599__A0 _03604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13323__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11610_ net1869 net1010 _07472_ _07475_ vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12590_ _03644_ net1843 net204 vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09464__B1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[5\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11271__B1 _07124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11541_ _07448_ _07451_ vssd1 vssd1 vccd1 vccd1 _07452_ sky130_fd_sc_hd__nor2_4
XFILLER_0_37_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_972 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14260_ net2936 _04019_ vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__nor2_1
X_11472_ net1001 _07382_ _07381_ vssd1 vssd1 vccd1 vccd1 _07383_ sky130_fd_sc_hd__a21oi_2
XANTENNA__09216__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13211_ _06536_ net2733 net353 vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__mux2_1
X_10423_ net896 _06439_ vssd1 vssd1 vccd1 vccd1 _06440_ sky130_fd_sc_hd__nor2_1
X_14191_ _07031_ net729 _03997_ _03998_ vssd1 vssd1 vccd1 vccd1 _00014_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_115_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11574__A1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13142_ net260 net2326 net447 vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__mux2_1
XANTENNA_input63_A wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10354_ _05982_ net510 _06125_ _06355_ _06373_ vssd1 vssd1 vccd1 vccd1 _06374_ sky130_fd_sc_hd__o221a_1
XFILLER_0_131_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17950_ clknet_leaf_35_wb_clk_i _03289_ _01646_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08990__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13073_ net254 net2411 net452 vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__mux2_1
X_10285_ _06197_ _06307_ net528 vssd1 vssd1 vccd1 vccd1 _06308_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_163_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12024_ _07834_ _07835_ vssd1 vssd1 vccd1 vccd1 _07836_ sky130_fd_sc_hd__or2_4
X_16901_ clknet_leaf_180_wb_clk_i _02531_ _00597_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_163_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_168_Right_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17881_ clknet_leaf_99_wb_clk_i _03224_ _01577_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08742__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10270__X _06294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_137_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16832_ clknet_leaf_131_wb_clk_i _02462_ _00528_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12402__S net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout590 _04368_ vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__buf_8
X_16763_ clknet_leaf_191_wb_clk_i _02393_ _00459_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13975_ _03845_ _03846_ vssd1 vssd1 vccd1 vccd1 _03847_ sky130_fd_sc_hd__nor2_1
X_15714_ net1152 vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12926_ net307 net2916 net473 vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__mux2_1
X_16694_ clknet_leaf_139_wb_clk_i _02324_ _00390_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13741__B _06609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15645_ net1248 vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__inv_2
X_12857_ net309 net2691 net480 vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__mux2_1
XANTENNA__13233__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18364_ net1349 vssd1 vssd1 vccd1 vccd1 la_data_out[12] sky130_fd_sc_hd__buf_2
XFILLER_0_56_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11808_ _07607_ _07609_ _07602_ vssd1 vssd1 vccd1 vccd1 _07620_ sky130_fd_sc_hd__a21oi_2
X_15576_ net1248 vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__inv_2
X_12788_ net330 net2595 net490 vssd1 vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__mux2_1
XANTENNA__12357__B _03650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10429__Y _06445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11262__B1 _07099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17315_ clknet_leaf_193_wb_clk_i _02945_ _01011_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_7_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11739_ _07542_ _07547_ _07550_ vssd1 vssd1 vccd1 vccd1 _07551_ sky130_fd_sc_hd__a21oi_1
X_14527_ net1182 vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18295_ net1387 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
XFILLER_0_43_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17246_ clknet_leaf_184_wb_clk_i _02876_ _00942_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14458_ net1052 vssd1 vssd1 vccd1 vccd1 _00088_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17586__D team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[23\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11014__B1 _06898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13409_ net2167 net260 net417 vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14389_ net1505 vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10445__X _06461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17177_ clknet_leaf_9_wb_clk_i _02807_ _00873_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11565__A1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16128_ net1306 vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_176_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08156__C_N team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08981__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08950_ _04990_ _05011_ vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__and2_1
X_16059_ net1262 vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12514__A0 _07789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08881_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[17\]
+ net801 net738 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_135_Right_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_102_Left_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13408__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08733__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire523_X net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09502_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[4\]
+ net673 net634 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[4\]
+ _05540_ vssd1 vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09433_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[5\]
+ net627 net609 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[5\]
+ _05475_ vssd1 vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13143__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09364_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[7\]
+ net811 net799 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05410_ sky130_fd_sc_hd__a22o_1
XANTENNA__09446__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_111_Left_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08315_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[31\]
+ net796 net791 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__a22o_1
XANTENNA__11253__B1 _07118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12982__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09295_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[8\]
+ net641 net600 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1257_A net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08246_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[31\]
+ net706 net697 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11005__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09576__B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08177_ _04252_ _04256_ net557 vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1045_X net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout884_A net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput160 net160 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__clkbuf_4
Xoutput171 net171 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_120_Left_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput182 net182 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10070_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[23\] _06098_ vssd1
+ vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout672_X net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13826__B net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13318__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08724__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09742__D net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10250__B _06273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout937_X net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13760_ _05212_ _06219_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[28\]
+ sky130_fd_sc_hd__and2_1
X_10972_ net1042 _06477_ _06953_ _06954_ vssd1 vssd1 vccd1 vccd1 _06955_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_69_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12711_ net283 net2646 net499 vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13691_ net1614 net1048 team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.next_state\[2\]
+ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_139_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13053__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12642_ net1690 _07836_ _03682_ vssd1 vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__mux2_1
X_15430_ net1124 vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15361_ net1228 vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_156_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12573_ _03650_ net1895 net206 vssd1 vssd1 vccd1 vccd1 _03068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12892__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17100_ clknet_leaf_5_wb_clk_i _02730_ _00796_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11524_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[26\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[26\]
+ net1033 vssd1 vssd1 vccd1 vccd1 _07435_ sky130_fd_sc_hd__mux2_1
X_14312_ _04083_ _04084_ vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18080_ clknet_leaf_83_wb_clk_i _00007_ _01776_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15292_ net1064 vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14243_ net2099 _04025_ vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__nor2_1
X_17031_ clknet_leaf_200_wb_clk_i _02661_ _00727_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11455_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[2\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[2\]
+ net1035 vssd1 vssd1 vccd1 vccd1 _07366_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10406_ net2866 net252 net539 vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__mux2_1
X_14174_ team_05_WB.instance_to_wrap.CPU_DAT_O\[23\] net504 net908 vssd1 vssd1 vccd1
+ vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[23\] sky130_fd_sc_hd__and3_1
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11386_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[9\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[8\]
+ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[4\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[7\]
+ vssd1 vssd1 vccd1 vccd1 _07317_ sky130_fd_sc_hd__or4b_1
XFILLER_0_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13125_ net326 net2441 net449 vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08963__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10337_ _06306_ _06357_ net521 vssd1 vssd1 vccd1 vccd1 _06358_ sky130_fd_sc_hd__mux2_1
X_17933_ clknet_leaf_43_wb_clk_i _03272_ _01629_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13056_ net331 net2249 net458 vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__mux2_1
X_10268_ net895 _06291_ vssd1 vssd1 vccd1 vccd1 _06292_ sky130_fd_sc_hd__nor2_1
XANTENNA__17492__Q team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[27\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12007_ net501 _07752_ _07770_ _07817_ _07818_ vssd1 vssd1 vccd1 vccd1 _07819_ sky130_fd_sc_hd__a221o_1
XANTENNA__08715__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13228__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11537__A _07379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17864_ clknet_leaf_104_wb_clk_i _03207_ _01560_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[46\]
+ sky130_fd_sc_hd__dfrtp_1
X_10199_ _06224_ vssd1 vssd1 vccd1 vccd1 _06225_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_159_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_159_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09652__D net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16815_ clknet_leaf_138_wb_clk_i _02445_ _00511_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_17795_ clknet_leaf_78_wb_clk_i _03138_ _01491_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[105\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_128_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13752__A _05212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16746_ clknet_leaf_17_wb_clk_i _02376_ _00442_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13958_ _04160_ _03830_ vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__nor2_1
XANTENNA__09140__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12909_ net261 net2581 net473 vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16677_ clknet_leaf_19_wb_clk_i _02307_ _00373_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13889_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[16\]
+ net558 net574 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[16\]
+ net985 vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__a221o_1
XANTENNA__14286__C _06408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15628_ net1150 vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09428__B1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11235__B1 _07125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18347_ net36 vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15559_ net1125 vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08100_ net1029 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[11\]
+ net976 _04199_ vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09080_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[13\]
+ net751 _04417_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__a22o_1
X_18278_ clknet_leaf_46_wb_clk_i _03507_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.key_data
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08031_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[18\] vssd1
+ vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__inv_2
Xinput40 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17229_ clknet_leaf_159_wb_clk_i _02859_ _00925_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput51 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
Xinput62 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold802 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2216 sky130_fd_sc_hd__dlygate4sd3_1
Xinput73 wbs_stb_i vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold813 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2227 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold824 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold835 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net2249 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold846 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2260 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10746__C1 _05924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold857 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 net2271 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08954__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold868 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net2282 sky130_fd_sc_hd__dlygate4sd3_1
X_09982_ _05442_ net361 vssd1 vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__nand2_1
Xhold879 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 net2293 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08933_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[16\]
+ net849 net798 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[16\]
+ _04994_ vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__a221o_1
XANTENNA__13138__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout298_A _06621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08706__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08864_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[17\]
+ net659 net633 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[17\]
+ _04928_ vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__a221o_1
Xhold1502 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 net2916 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1513 net76 vssd1 vssd1 vccd1 vccd1 net2927 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1524 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 net2938 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1535 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2949 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1546 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 net2960 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1557 team_05_WB.instance_to_wrap.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 net2971
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08795_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[19\]
+ net798 net741 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[19\]
+ _04864_ vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__a221o_1
XANTENNA__12977__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout465_A _03710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09667__B1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_2_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout632_A net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09416_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[6\]
+ net814 net791 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[6\]
+ _05459_ vssd1 vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08194__C team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[25\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11226__B1 _07126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09347_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[7\]
+ net669 _05393_ net721 vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__a211o_1
XANTENNA__09858__Y _05887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout420_X net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13601__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08642__A1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09278_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[9\]
+ net797 _05325_ _05327_ net855 vssd1 vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_62_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08229_ net887 net866 _04294_ vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_151_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11240_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[52\] _07110_
+ _07124_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[28\] _07202_
+ vssd1 vssd1 vccd1 vccd1 _07203_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09198__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08945__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11171_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[55\] _07117_
+ _07120_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[39\] vssd1 vssd1
+ vccd1 vccd1 _07137_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10122_ _04818_ net364 vssd1 vssd1 vccd1 vccd1 _06150_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09753__C net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13048__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14930_ net1233 vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__inv_2
X_10053_ _06047_ net337 _06066_ _06081_ vssd1 vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__o211a_1
XANTENNA__11701__A1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[31\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input26_A DAT_I[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09370__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14861_ net1080 vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__inv_2
XANTENNA__12887__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16600_ clknet_leaf_27_wb_clk_i _02230_ _00296_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13812_ net1594 net971 net724 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[23\]
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_106_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17580_ clknet_leaf_72_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[17\]
+ _01276_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14792_ net1224 vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16531_ clknet_leaf_165_wb_clk_i _02161_ _00227_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09122__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13743_ net922 _06572_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[11\]
+ sky130_fd_sc_hd__nor2_1
X_10955_ net1042 _06420_ vssd1 vssd1 vccd1 vccd1 _06941_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_27_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_158_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_123_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12009__A2 _07623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16462_ clknet_leaf_171_wb_clk_i _02092_ _00158_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10886_ _06783_ _06882_ _06781_ vssd1 vssd1 vccd1 vccd1 _06883_ sky130_fd_sc_hd__o21ai_1
X_13674_ net2097 net269 net384 vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18201_ clknet_leaf_33_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[22\]
+ _01896_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_15413_ net1138 vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__inv_2
XANTENNA__11217__B1 _07104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12625_ _03620_ net1864 net201 vssd1 vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12475__X _03674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16393_ clknet_leaf_20_wb_clk_i _02023_ _00089_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13511__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18132_ clknet_leaf_48_wb_clk_i _00028_ _01828_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12556_ _03644_ net1771 net205 vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__mux2_1
X_15344_ net1183 vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09830__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11507_ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[12\] _07417_ net1001
+ vssd1 vssd1 vccd1 vccd1 _07418_ sky130_fd_sc_hd__mux2_1
XANTENNA__10440__A1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18063_ clknet_leaf_86_wb_clk_i _03401_ _01759_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__dfrtp_1
X_12487_ net2098 _03644_ net211 vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15275_ net1076 vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__inv_2
XANTENNA__09647__D net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold109 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1523 sky130_fd_sc_hd__dlygate4sd3_1
X_17014_ clknet_leaf_143_wb_clk_i _02644_ _00710_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09189__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14226_ team_05_WB.instance_to_wrap.total_design.keypad0.counter\[9\] _04021_ vssd1
+ vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__and2_1
X_11438_ net1050 net1049 team_05_WB.instance_to_wrap.total_design.core.instr_fetch
+ vssd1 vssd1 vccd1 vccd1 _07351_ sky130_fd_sc_hd__or3_4
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08397__B1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13747__A net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14157_ _03910_ _03994_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[6\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__08936__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11369_ net957 _06743_ _07307_ vssd1 vssd1 vccd1 vccd1 _07308_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13108_ net264 net2522 net448 vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__mux2_1
X_14088_ _03938_ _03952_ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__nor2_1
X_17916_ clknet_leaf_51_wb_clk_i _00000_ _01612_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.wishbone.curr_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_13039_ net246 net2893 net458 vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13693__A1 team_05_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1160 net1161 vssd1 vssd1 vccd1 vccd1 net1160 sky130_fd_sc_hd__buf_4
Xfanout1171 net1174 vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__buf_4
XANTENNA__09361__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17847_ clknet_leaf_89_wb_clk_i _03190_ _01543_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[93\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1182 net1186 vssd1 vssd1 vccd1 vccd1 net1182 sky130_fd_sc_hd__buf_4
XANTENNA__12797__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1193 net1194 vssd1 vssd1 vccd1 vccd1 net1193 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11554__X _07465_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08580_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[25\]
+ net717 _04646_ _04655_ vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__o22ai_4
X_17778_ clknet_leaf_95_wb_clk_i _03121_ _01474_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12369__Y _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14297__B team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[31\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09113__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16729_ clknet_leaf_9_wb_clk_i _02359_ _00425_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08295__B net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09201_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[10\]
+ net683 _05253_ net720 vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__a211o_1
XANTENNA__11208__B1 _07106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_56_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_146_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13421__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09132_ _05165_ _05185_ vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__and2_1
XFILLER_0_127_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09821__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10617__Y _06623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09063_ _05118_ _05119_ _05120_ _05121_ vssd1 vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__or4_1
XFILLER_0_163_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout213_A _03671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold610 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2024 sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2035 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold632 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2046 sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net2057 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13920__A2 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold654 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2068 sky130_fd_sc_hd__dlygate4sd3_1
Xhold665 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2079 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold676 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2090 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1122_A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold687 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 net2101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold698 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2112 sky130_fd_sc_hd__dlygate4sd3_1
X_09965_ _05909_ _05993_ vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout582_A _03761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08916_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[16\]
+ net707 net660 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[16\]
+ _04980_ vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__a221o_1
X_09896_ _04273_ _05923_ vssd1 vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__nand2_1
Xhold1310 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net2724 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1321 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 net2735 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10498__B2 _06060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1332 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net2746 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1343 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2757 sky130_fd_sc_hd__dlygate4sd3_1
X_08847_ _04908_ _04910_ _04912_ _04914_ vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__or4_1
Xhold1354 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 net2768 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14488__A net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout847_A _04373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout468_X net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1365 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2779 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1376 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2790 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12500__S _03674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08778_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[19\]
+ net704 net632 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[19\]
+ _04848_ vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__a221o_1
Xhold1387 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2801 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1398 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2812 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09104__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18403__1373 vssd1 vssd1 vccd1 vccd1 _18403__1373/HI net1373 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_0_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout635_X net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_3_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_0_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11998__A1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[17\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10740_ net1018 _05733_ net551 vssd1 vssd1 vccd1 vccd1 _06739_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10671_ _05951_ _06673_ net894 vssd1 vssd1 vccd1 vccd1 _06674_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout802_X net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12410_ net1680 _07789_ _03667_ vssd1 vssd1 vccd1 vccd1 _03220_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13331__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13390_ net2202 net311 net420 vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09812__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09748__C _04287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12341_ _03536_ _03540_ _03530_ vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15060_ net1073 vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12272_ _03559_ _03566_ vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14011_ _03860_ _03881_ vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__nand2_1
XANTENNA__08379__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11223_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[77\] _07116_
+ _07121_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[85\] _07186_
+ vssd1 vssd1 vccd1 vccd1 _07187_ sky130_fd_sc_hd__a221o_1
XANTENNA__08918__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10543__X _06554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10186__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11154_ _07080_ _07112_ vssd1 vssd1 vccd1 vccd1 _07120_ sky130_fd_sc_hd__nor2_4
XANTENNA__09591__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10105_ _05078_ net364 vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__or2_1
X_11085_ _07040_ _07042_ _07051_ _04161_ vssd1 vssd1 vccd1 vccd1 _07052_ sky130_fd_sc_hd__a2bb2o_2
X_15962_ net1289 vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17701_ clknet_leaf_101_wb_clk_i _03044_ _01397_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09780__A _05442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10036_ net371 _06062_ vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__nand2_1
XANTENNA__09343__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14913_ net1219 vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__inv_2
X_15893_ net1295 vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_125_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13506__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08551__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17632_ clknet_leaf_54_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.branch_ff
+ _01328_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.program_count.ALU_out_reg
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12410__S _03667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14844_ net1083 vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17563_ clknet_leaf_115_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[0\]
+ _01259_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14775_ net1102 vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11987_ _07777_ _07785_ _07795_ vssd1 vssd1 vccd1 vccd1 _07799_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08303__B1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11989__A1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[21\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16514_ clknet_leaf_6_wb_clk_i _02144_ _00210_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13726_ net906 _06273_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[26\]
+ sky130_fd_sc_hd__and2_1
X_10938_ net956 _06350_ vssd1 vssd1 vccd1 vccd1 _06927_ sky130_fd_sc_hd__nor2_1
XANTENNA__08854__A1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17494_ clknet_leaf_37_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[29\]
+ _01190_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_79 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16445_ clknet_leaf_131_wb_clk_i _02075_ _00141_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10869_ _06809_ _06865_ _06806_ _06807_ vssd1 vssd1 vccd1 vccd1 _06866_ sky130_fd_sc_hd__o211a_1
XFILLER_0_112_1053 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13657_ net2890 net307 net389 vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__mux2_1
XANTENNA__09899__A_N _04613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13241__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12608_ net1727 _07836_ _03680_ vssd1 vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_951 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16376_ clknet_leaf_27_wb_clk_i _02006_ _00072_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13588_ net2187 net310 net396 vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18115_ clknet_leaf_45_wb_clk_i _00005_ _01811_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.key_confirm
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11610__B1 _07472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15327_ net1180 vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__inv_2
X_12539_ _07836_ net1870 _03675_ vssd1 vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__mux2_1
XANTENNA__08082__A2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[20\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18046_ net1039 _03384_ _01742_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_124_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15258_ net1053 vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17594__D team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[31\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14209_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[10\] _04008_
+ _04009_ vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__o21a_1
XANTENNA__08909__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13902__A2 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09674__B net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15189_ net1059 vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_174_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_174_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout408 _03728_ vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__buf_8
XANTENNA__08153__A_N net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout419 _03726_ vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_103_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_103_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08790__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09750_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[0\]
+ net886 net875 net870 vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__and4_1
XANTENNA__09334__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08701_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[22\]
+ net661 net604 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[22\]
+ _04762_ vssd1 vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_33_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09681_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[1\]
+ net878 net872 net858 vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__and4_1
XANTENNA__08542__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11725__A _07379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08632_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[24\]
+ net799 net766 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[24\]
+ _04703_ vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__a221o_1
XANTENNA__13416__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08563_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[25\]
+ net705 net662 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[25\]
+ _04638_ vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_81_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08494_ _04559_ _04560_ _04570_ _04571_ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__or4_2
XFILLER_0_162_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout330_A _06705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout428_A net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13151__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1072_A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09568__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09115_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[12\]
+ net771 net741 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[12\]
+ _05167_ vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__a221o_1
XANTENNA__11601__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12990__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10076__A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14771__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout216_X net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09046_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[13\]
+ net632 net614 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout797_A _04395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold440 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[39\] vssd1 vssd1
+ vccd1 vccd1 net1854 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09584__B net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold451 team_05_WB.instance_to_wrap.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 net1865
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13818__C net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold462 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1876 sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 net162 vssd1 vssd1 vccd1 vccd1 net1887 sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[125\] vssd1 vssd1
+ vccd1 vccd1 net1898 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold495 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[5\] vssd1 vssd1
+ vccd1 vccd1 net1909 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout920 _07352_ vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__buf_2
Xfanout931 _04374_ vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08781__B1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09948_ _05930_ _05974_ _05884_ _05887_ vssd1 vssd1 vccd1 vccd1 _05977_ sky130_fd_sc_hd__o211a_1
Xfanout942 net943 vssd1 vssd1 vccd1 vccd1 net942 sky130_fd_sc_hd__clkbuf_2
Xfanout953 net955 vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__buf_2
XANTENNA__13657__A1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout964 _04243_ vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__buf_2
Xfanout975 net977 vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__buf_2
Xfanout986 net987 vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_146_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09879_ _04634_ _05907_ vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__nor2_1
Xfanout997 net999 vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout752_X net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1140 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2554 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08533__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11635__A team_05_WB.instance_to_wrap.wishbone.curr_state\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1151 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2565 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13326__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11910_ _07529_ _07721_ vssd1 vssd1 vccd1 vccd1 _07722_ sky130_fd_sc_hd__nor2_1
Xhold1162 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 net2576 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1173 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 net2587 sky130_fd_sc_hd__dlygate4sd3_1
X_12890_ net311 net2354 net476 vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1184 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2598 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09750__D net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1195 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 net2609 sky130_fd_sc_hd__dlygate4sd3_1
X_11841_ _07620_ _07624_ _07628_ _07623_ vssd1 vssd1 vccd1 vccd1 _07653_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_16_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09599__X _05634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14560_ net1102 vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__inv_2
X_11772_ _07569_ _07571_ _07565_ vssd1 vssd1 vccd1 vccd1 _07584_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13511_ net2558 net274 net406 vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__mux2_1
X_10723_ _06112_ _06121_ vssd1 vssd1 vccd1 vccd1 _06723_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14491_ net1095 vssd1 vssd1 vccd1 vccd1 _00121_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16230_ net1202 vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__inv_2
X_10654_ _05809_ _05813_ vssd1 vssd1 vccd1 vccd1 _06658_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_125_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13442_ net2801 net259 net412 vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__mux2_1
XANTENNA__11199__A2 _07117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12396__B2 _07914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16161_ net1164 vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__inv_2
X_13373_ net2675 net254 net420 vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__mux2_1
X_10585_ net892 _06590_ _06592_ vssd1 vssd1 vccd1 vccd1 _06593_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload18 clknet_leaf_203_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload18/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__10946__A2 _06369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload29 clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload29/Y sky130_fd_sc_hd__inv_8
X_15112_ net1218 vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__inv_2
X_12324_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[19\] net1000 _03588_
+ net543 vssd1 vssd1 vccd1 vccd1 _03619_ sky130_fd_sc_hd__a211oi_2
XTAP_TAPCELL_ROW_118_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16092_ net1308 vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_1_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_51_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12255_ _03516_ _03537_ _03547_ _03549_ vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__nor4_1
XFILLER_0_121_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15043_ net1204 vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_43_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_50_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11206_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[5\] _07092_ _07124_
+ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[29\] vssd1 vssd1 vccd1
+ vccd1 _07170_ sky130_fd_sc_hd__a22o_1
X_12186_ _07936_ _07940_ _07996_ vssd1 vssd1 vccd1 vccd1 _07998_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08772__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11137_ _07059_ _07068_ _07071_ vssd1 vssd1 vccd1 vccd1 _07103_ sky130_fd_sc_hd__and3_4
X_16994_ clknet_leaf_5_wb_clk_i _02624_ _00690_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09316__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11068_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[2\] _07034_
+ vssd1 vssd1 vccd1 vccd1 _07035_ sky130_fd_sc_hd__or2_2
X_15945_ net1266 vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__inv_2
XANTENNA__11123__A2 _07031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13236__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08524__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11545__A net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10019_ _05531_ _06002_ vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__nor2_1
XANTENNA__15017__A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15876_ net1293 vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__inv_2
X_17615_ clknet_leaf_49_wb_clk_i _02986_ _01311_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_14827_ net1067 vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__inv_2
XANTENNA__13760__A _05212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17546_ clknet_leaf_49_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[17\]
+ _01242_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_148_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14758_ net1247 vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17589__D team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[26\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13709_ net901 _06609_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[9\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17477_ clknet_leaf_39_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[12\]
+ _01173_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14689_ net1223 vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16428_ clknet_leaf_2_wb_clk_i _02058_ _00124_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_82_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_73_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12387__A1 _03663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16359_ clknet_leaf_200_wb_clk_i _01989_ _00055_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18029_ clknet_leaf_97_wb_clk_i _03368_ _01725_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout205 net207 vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__clkbuf_4
Xfanout216 net217 vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__buf_4
XANTENNA__08763__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09802_ _05146_ _05830_ vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__nor2_2
Xfanout227 net229 vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout238 net241 vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__clkbuf_2
Xfanout249 _06405_ vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10570__B1 _06051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09733_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[0\]
+ net836 net771 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_2_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13146__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09664_ net588 _05695_ _05696_ _05697_ vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__nand4_1
XANTENNA__09570__D net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08615_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[24\]
+ net701 net638 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[24\]
+ _04689_ vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__a221o_1
XANTENNA__12985__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09595_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[2\]
+ net826 _05605_ _05609_ _05618_ vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__a2111o_1
Xclkbuf_leaf_71_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout545_A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1287_A net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08546_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[26\]
+ net743 net740 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08477_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[27\]
+ net669 net622 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__a22o_1
XANTENNA__09579__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout333_X net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout712_A _04288_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12378__A1 _03610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout500_X net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11050__A1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_149_Right_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10370_ net888 _05977_ _05978_ _06388_ vssd1 vssd1 vccd1 vccd1 _06389_ sky130_fd_sc_hd__or4_1
XANTENNA__13829__B net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09029_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[14\]
+ net783 net761 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_148_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09745__D net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12040_ net919 _07849_ _07850_ _07840_ _07847_ vssd1 vssd1 vccd1 vccd1 _07852_ sky130_fd_sc_hd__o2111a_4
XTAP_TAPCELL_ROW_148_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold270 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[114\] vssd1 vssd1
+ vccd1 vccd1 net1684 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09546__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold281 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[0\] vssd1 vssd1
+ vccd1 vccd1 net1695 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[117\] vssd1 vssd1
+ vccd1 vccd1 net1706 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_72_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12550__A1 _07791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08754__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_127_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout750 net751 vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__clkbuf_4
Xfanout761 net763 vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__clkbuf_8
Xfanout772 _04406_ vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__clkbuf_8
X_13991_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[6\] _03840_ _03861_
+ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__o21a_1
Xfanout783 net785 vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__buf_6
XFILLER_0_99_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout794 net795 vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08506__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13056__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15730_ net1295 vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_161_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12942_ net255 net2611 net468 vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_161_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15661_ net1140 vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12895__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12873_ net253 net2459 net476 vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__mux2_1
X_17400_ clknet_leaf_56_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[0\]
+ _01096_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14612_ net1075 vssd1 vssd1 vccd1 vccd1 _00242_ sky130_fd_sc_hd__inv_2
XANTENNA__08809__A1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18380_ net1365 vssd1 vssd1 vccd1 vccd1 la_data_out[28] sky130_fd_sc_hd__buf_2
X_11824_ _07633_ _07634_ _07619_ vssd1 vssd1 vccd1 vccd1 _07636_ sky130_fd_sc_hd__a21o_1
X_15592_ net1245 vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17331_ clknet_leaf_169_wb_clk_i _02961_ _01027_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[27\]
+ sky130_fd_sc_hd__dfrtp_2
X_14543_ net1286 vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__inv_2
XANTENNA__08285__A2 _04347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11755_ _07565_ _07566_ vssd1 vssd1 vccd1 vccd1 _07567_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17262_ clknet_leaf_177_wb_clk_i _02892_ _00958_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14358__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10706_ _05806_ _05948_ vssd1 vssd1 vccd1 vccd1 _06707_ sky130_fd_sc_hd__xnor2_1
X_14474_ net1111 vssd1 vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__inv_2
X_11686_ net47 net49 net48 net46 vssd1 vssd1 vccd1 vccd1 _07500_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_24_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16213_ net1085 vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13425_ net2755 net325 net417 vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10637_ net890 _06641_ _06640_ net555 vssd1 vssd1 vccd1 vccd1 _06642_ sky130_fd_sc_hd__a211o_1
X_17193_ clknet_leaf_25_wb_clk_i _02823_ _00889_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload107 clknet_leaf_159_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload107/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__10919__A2 _06907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload118 clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload118/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_23_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16144_ net1273 vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__inv_2
Xclkload129 clknet_leaf_139_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload129/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_107_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10568_ _06049_ _06254_ vssd1 vssd1 vccd1 vccd1 _06577_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13356_ net328 net2912 net426 vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_166_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12307_ _03590_ _03601_ vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16075_ net1173 vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10499_ _06359_ _06503_ _06506_ net335 _06511_ vssd1 vssd1 vccd1 vccd1 _06512_ sky130_fd_sc_hd__o221a_1
X_13287_ net303 net2606 net434 vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_15_Left_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09537__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15026_ net1238 vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__inv_2
X_12238_ _03519_ _03524_ _03527_ vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__and3_1
XANTENNA__12541__A1 _03623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13755__A _05212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12169_ _07979_ _07980_ vssd1 vssd1 vccd1 vccd1 _07981_ sky130_fd_sc_hd__nor2_1
XANTENNA__10552__B1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16977_ clknet_leaf_123_wb_clk_i _02607_ _00673_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09671__C net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14289__C _06108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput5 DAT_I[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
X_15928_ net1266 vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__inv_2
XANTENNA__09170__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15859_ net1303 vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__inv_2
XANTENNA__14586__A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08400_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[29\]
+ net663 net637 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__a22o_1
X_09380_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[6\]
+ net707 net630 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05425_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08331_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[31\]
+ net762 net757 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17529_ clknet_leaf_60_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[0\]
+ _01225_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_7_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08262_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[31\] _04269_
+ vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__and2_2
XANTENNA__10083__A2 _06108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08193_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[13\] _04274_
+ _04239_ vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16306__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10057__C team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11032__A1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08984__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1035_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09565__D net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09528__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08736__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout495_A _03699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09862__B _05888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08200__A2 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16041__A net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1202_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09207__X _05260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09581__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout283_X net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout662_A net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09716_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[0\]
+ net950 net939 net931 vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__and4_1
XFILLER_0_69_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09647_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[1\]
+ net1015 net946 net927 vssd1 vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout450_X net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout927_A net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13604__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09578_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[2\]
+ net1015 net946 net932 vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__and4_1
XFILLER_0_93_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08529_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[26\]
+ net670 net639 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[26\]
+ _04605_ vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09464__A1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout715_X net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11540_ _07380_ _07450_ vssd1 vssd1 vccd1 vccd1 _07451_ sky130_fd_sc_hd__nor2_8
XFILLER_0_9_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11471_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[0\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[0\]
+ net1033 vssd1 vssd1 vccd1 vccd1 _07382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10422_ _06096_ _06438_ vssd1 vssd1 vccd1 vccd1 _06439_ sky130_fd_sc_hd__or2_1
X_13210_ net272 net2516 net350 vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09767__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14190_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[3\] _07027_
+ vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_115_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11574__A2 _07354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08975__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10353_ _06051_ _06372_ vssd1 vssd1 vccd1 vccd1 _06373_ sky130_fd_sc_hd__nand2_1
X_13141_ net265 net2904 net447 vssd1 vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_111_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09519__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13072_ net248 net2488 net454 vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__mux2_1
XANTENNA_input56_A wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10284_ _06259_ _06306_ net521 vssd1 vssd1 vccd1 vccd1 _06307_ sky130_fd_sc_hd__mux2_1
XANTENNA__12523__A1 _03614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12023_ net356 _07736_ vssd1 vssd1 vccd1 vccd1 _07835_ sky130_fd_sc_hd__nor2_1
X_16900_ clknet_leaf_194_wb_clk_i _02530_ _00596_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17880_ clknet_leaf_92_wb_clk_i _03223_ _01576_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_163_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16831_ clknet_leaf_153_wb_clk_i _02461_ _00527_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout580 net581 vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__clkbuf_2
Xfanout591 _04368_ vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__clkbuf_4
X_16762_ clknet_leaf_10_wb_clk_i _02392_ _00458_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13974_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[10\] _03844_ vssd1
+ vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__nor2_1
X_15713_ net1153 vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__inv_2
X_12925_ net326 net2406 net473 vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1091 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16693_ clknet_leaf_71_wb_clk_i _02323_ _00389_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13514__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15644_ net1248 vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__inv_2
X_12856_ net329 net2778 net482 vssd1 vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18363_ net1348 vssd1 vssd1 vccd1 vccd1 la_data_out[11] sky130_fd_sc_hd__buf_2
X_11807_ _07614_ _07618_ _07615_ vssd1 vssd1 vccd1 vccd1 _07619_ sky130_fd_sc_hd__o21a_1
XFILLER_0_150_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15575_ net1251 vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12787_ net315 net2762 net491 vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12357__C _03651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17314_ clknet_leaf_15_wb_clk_i _02944_ _01010_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14526_ net1068 vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11738_ _07532_ _07549_ _07542_ vssd1 vssd1 vccd1 vccd1 _07550_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_25_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18294_ net1386 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
XFILLER_0_25_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17245_ clknet_leaf_128_wb_clk_i _02875_ _00941_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09207__A1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[30\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14457_ net1051 vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12654__A _07346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11669_ net2 net989 net916 net1890 vssd1 vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__o22a_1
XFILLER_0_126_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13408_ net2296 net265 net416 vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17176_ clknet_leaf_29_wb_clk_i _02806_ _00872_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14388_ net1521 vssd1 vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11565__A2 _07354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08966__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16127_ net1307 vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__inv_2
X_13339_ net248 net2373 net426 vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__mux2_1
XANTENNA__08430__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16058_ net1262 vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__inv_2
XANTENNA__17953__Q net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11317__A2 _07106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08718__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11557__X _07468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15009_ net1235 vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__inv_2
X_08880_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[29\] net965
+ net955 _04946_ _04345_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[17\]
+ sky130_fd_sc_hd__a221o_1
XANTENNA_wire349_X net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_74 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10113__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09143__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09501_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[4\]
+ net708 net657 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__a22o_1
XANTENNA__12388__X _03664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08497__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13424__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09432_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[5\]
+ net705 net612 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05475_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09363_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[7\]
+ net783 net765 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[7\]
+ _05408_ vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08249__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08314_ net1016 net949 net933 vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_23_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09294_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[8\]
+ net612 net609 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[8\]
+ _05342_ vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__a221o_1
XANTENNA_10 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08245_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[31\]
+ net649 net595 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[31\]
+ _04327_ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout410_A _03728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1152_A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16036__A net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11005__A1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08406__C1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08176_ team_05_WB.instance_to_wrap.total_design.core.instr_fetch _04258_ vssd1 vssd1
+ vccd1 vccd1 _04259_ sky130_fd_sc_hd__nor2_1
XFILLER_0_144_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09576__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08957__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08421__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10084__A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09873__A _04656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput150 net150 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
Xoutput161 net161 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
XANTENNA__11308__A2 _07100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12505__A1 _07836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08709__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout877_A net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput172 net172 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout498_X net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput183 net914 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__clkbuf_4
XANTENNA__12503__S _03673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10371__X _06390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09382__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09921__A2 _05949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout665_X net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10971_ _06804_ _06805_ _06867_ net1042 vssd1 vssd1 vccd1 vccd1 _06954_ sky130_fd_sc_hd__o31a_1
XANTENNA__08488__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout832_X net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08495__Y _04573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13334__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12710_ net274 net2888 net498 vssd1 vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13690_ net2915 net307 net387 vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_139_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12641_ _03650_ net1709 net201 vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_139_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15360_ net1103 vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12572_ net1717 _07816_ _03678_ vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_156_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09400__X team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14311_ _04777_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[22\]
+ _04818_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__o22a_1
X_11523_ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[15\] _07433_ net1001
+ vssd1 vssd1 vccd1 vccd1 _07434_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15291_ net1099 vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__inv_2
XANTENNA__12474__A _07840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08660__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17030_ clknet_leaf_117_wb_clk_i _02660_ _00726_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14242_ _04021_ _04031_ vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__nor2_1
X_11454_ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[3\] _07364_ net1002
+ vssd1 vssd1 vccd1 vccd1 _07365_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08948__B1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[16\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10405_ net382 _06422_ vssd1 vssd1 vccd1 vccd1 _06423_ sky130_fd_sc_hd__and2_1
X_11385_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[17\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[16\]
+ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[15\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[14\]
+ vssd1 vssd1 vccd1 vccd1 _07316_ sky130_fd_sc_hd__or4_1
X_14173_ net1791 net502 net908 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[22\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__08412__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13124_ net321 net1979 net449 vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__mux2_1
X_10336_ _06041_ _06078_ vssd1 vssd1 vccd1 vccd1 _06357_ sky130_fd_sc_hd__nor2_1
XANTENNA__13509__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12413__S _03667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10267_ _06101_ _06290_ vssd1 vssd1 vccd1 vccd1 _06291_ sky130_fd_sc_hd__or2_1
X_17932_ clknet_leaf_43_wb_clk_i _03271_ _01628_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13055_ net313 net2861 net459 vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__mux2_1
X_12006_ _07765_ _07773_ vssd1 vssd1 vccd1 vccd1 _07818_ sky130_fd_sc_hd__nor2_1
X_17863_ clknet_leaf_88_wb_clk_i _03206_ _01559_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11537__B _07447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10198_ _06222_ _06223_ net526 vssd1 vssd1 vccd1 vccd1 _06224_ sky130_fd_sc_hd__mux2_1
XANTENNA__11180__B1 _07111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13592__X _03732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16814_ clknet_leaf_175_wb_clk_i _02444_ _00510_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_17794_ clknet_leaf_92_wb_clk_i _03137_ _01490_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[104\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09125__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13752__B _06408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16745_ clknet_leaf_14_wb_clk_i _02375_ _00441_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13957_ _03828_ _03829_ vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__or2_1
XANTENNA__08479__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13244__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11553__A _07348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_199_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_199_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12908_ net265 net2250 net472 vssd1 vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__mux2_1
X_16676_ clknet_leaf_183_wb_clk_i _02306_ _00372_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13888_ net1576 net982 _03780_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[15\]
+ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_128_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_128_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15627_ net1149 vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12839_ net247 net2796 net481 vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18346_ net35 vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15558_ net1116 vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17948__Q team_05_WB.instance_to_wrap.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14509_ net1087 vssd1 vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__inv_2
X_18277_ clknet_leaf_42_wb_clk_i _03506_ _01972_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[31\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09677__B net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15489_ net1154 vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__inv_2
XANTENNA__08651__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08030_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[19\] vssd1
+ vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17228_ clknet_leaf_2_wb_clk_i _02858_ _00924_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput30 DAT_I[6] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput41 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput52 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__buf_1
Xinput63 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08939__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold803 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net2217 sky130_fd_sc_hd__dlygate4sd3_1
Xinput74 wbs_we_i vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__buf_1
X_17159_ clknet_leaf_202_wb_clk_i _02789_ _00855_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold814 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 net2228 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold825 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2239 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08403__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold836 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net2261 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold858 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2272 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold869 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2283 sky130_fd_sc_hd__dlygate4sd3_1
X_09981_ net375 net365 vssd1 vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__nand2_1
XANTENNA__10903__Y _06898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13419__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08932_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[16\]
+ net778 net764 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[16\]
+ _04995_ vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__a221o_1
XANTENNA__10632__A _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09364__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08863_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[17\]
+ net665 net647 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[17\]
+ _04929_ vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__a221o_1
Xhold1503 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net2917 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11171__B1 _07120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout193_A _06184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1514 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 net2928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1525 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2939 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1536 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1547 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 net2961 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1558 team_05_WB.instance_to_wrap.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 net2972
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08794_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[19\]
+ net849 net802 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__a22o_1
XANTENNA__09116__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09667__A1 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11463__A net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout458_A _03712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13154__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11474__A1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09415_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[6\]
+ net775 net761 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__a22o_1
XANTENNA__12993__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout625_A net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08890__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09346_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[7\]
+ net618 net595 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_62_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09277_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[9\]
+ net766 net762 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[9\]
+ _05326_ vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout413_X net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08642__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[24\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08228_ net879 net869 net867 vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__and3_1
XFILLER_0_62_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout994_A _07470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08159_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[4\] team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[2\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[6\] team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__and4b_1
XFILLER_0_132_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11170_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[79\] _07116_
+ _07119_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[31\] _07135_
+ vssd1 vssd1 vccd1 vccd1 _07136_ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout782_X net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13329__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10121_ _04777_ net367 vssd1 vssd1 vccd1 vccd1 _06149_ sky130_fd_sc_hd__nand2_1
XFILLER_0_140_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09753__D _04296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09355__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10052_ net524 _06080_ net333 _06072_ vssd1 vssd1 vccd1 vccd1 _06081_ sky130_fd_sc_hd__a211o_1
XANTENNA__11701__A2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[25\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14860_ net1078 vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__inv_2
X_13811_ net1607 net970 net723 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[22\]
+ sky130_fd_sc_hd__and3_1
XANTENNA_input19_A DAT_I[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14791_ net1199 vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13064__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16530_ clknet_leaf_121_wb_clk_i _02160_ _00226_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13742_ net923 _06591_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[10\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_27_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10954_ _06799_ _06872_ vssd1 vssd1 vccd1 vccd1 _06940_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_27_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16461_ clknet_leaf_162_wb_clk_i _02091_ _00157_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13673_ net2236 net259 net387 vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__mux2_1
X_10885_ _06784_ _06880_ _06782_ vssd1 vssd1 vccd1 vccd1 _06882_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08881__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18200_ clknet_leaf_36_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[21\]
+ _01895_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_15412_ net1131 vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__inv_2
XANTENNA__12414__A0 _03646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12624_ _03644_ net1916 net202 vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16392_ clknet_leaf_203_wb_clk_i _02022_ _00088_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08618__C1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18131_ clknet_leaf_48_wb_clk_i _00027_ _01827_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15343_ net1233 vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__inv_2
X_12555_ _03610_ net1875 net205 vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12408__S net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10717__A team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08633__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11506_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[12\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[12\]
+ net1034 vssd1 vssd1 vccd1 vccd1 _07417_ sky130_fd_sc_hd__mux2_1
X_18062_ clknet_leaf_99_wb_clk_i _03400_ _01758_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15274_ net1121 vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12486_ net1706 _03610_ net211 vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__mux2_1
X_17013_ clknet_leaf_23_wb_clk_i _02643_ _00709_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_14225_ team_05_WB.instance_to_wrap.total_design.keypad0.counter\[7\] team_05_WB.instance_to_wrap.total_design.keypad0.counter\[8\]
+ _04020_ vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11437_ _07349_ vssd1 vssd1 vccd1 vccd1 _07350_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10728__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13747__B _06500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14156_ _03882_ _03994_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[5\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11368_ _06841_ _06899_ _07306_ vssd1 vssd1 vccd1 vccd1 _07307_ sky130_fd_sc_hd__or3b_1
XFILLER_0_42_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13107_ net255 net2159 net448 vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__mux2_1
XANTENNA__13239__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10319_ net556 _06323_ _06340_ vssd1 vssd1 vccd1 vccd1 _06341_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14087_ _03932_ _03950_ _03951_ vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__and3_1
X_11299_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[73\] _07116_
+ _07121_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[81\] _07258_
+ vssd1 vssd1 vccd1 vccd1 _07259_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09346__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17915_ clknet_leaf_63_wb_clk_i _00003_ _01611_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09018__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[14\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13038_ net228 net2567 net458 vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__mux2_1
Xfanout1150 net1151 vssd1 vssd1 vccd1 vccd1 net1150 sky130_fd_sc_hd__buf_2
XANTENNA__13693__A2 _00040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13763__A net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1161 net1162 vssd1 vssd1 vccd1 vccd1 net1161 sky130_fd_sc_hd__clkbuf_4
Xfanout1172 net1174 vssd1 vssd1 vccd1 vccd1 net1172 sky130_fd_sc_hd__clkbuf_4
X_17846_ clknet_leaf_74_wb_clk_i _03189_ _01542_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[92\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08857__A net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1183 net1186 vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__clkbuf_4
Xfanout1194 net1211 vssd1 vssd1 vccd1 vccd1 net1194 sky130_fd_sc_hd__clkbuf_4
X_17777_ clknet_leaf_99_wb_clk_i _03120_ _01473_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_14989_ net1082 vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16728_ clknet_leaf_28_wb_clk_i _02358_ _00424_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16659_ clknet_leaf_164_wb_clk_i _02289_ _00355_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09200_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[10\]
+ net691 net605 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09131_ _05165_ _05185_ vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_40_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18329_ team_05_WB.instance_to_wrap.lcd_en vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08624__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09062_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[13\]
+ net660 net624 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[13\]
+ _05106_ vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__a221o_1
XFILLER_0_142_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_96_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_7_Left_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold600 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2014 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout206_A net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10719__B1 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold611 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net2025 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_25_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_114_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold622 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net2036 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold633 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net2047 sky130_fd_sc_hd__dlygate4sd3_1
Xhold644 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[79\] vssd1 vssd1
+ vccd1 vccd1 net2058 sky130_fd_sc_hd__dlygate4sd3_1
Xhold655 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net2069 sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2080 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13149__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold677 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 net2091 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold688 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 net2102 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09964_ _04573_ _04592_ _05992_ vssd1 vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__a21bo_1
Xhold699 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 net2113 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09573__D net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09337__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08915_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[16\]
+ net664 net640 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__a22o_1
X_09895_ _04273_ _05923_ vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__and2_4
XANTENNA__12988__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1300 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 net2714 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1311 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 net2725 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1322 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net2736 sky130_fd_sc_hd__dlygate4sd3_1
X_08846_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[18\]
+ net841 net786 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[18\]
+ _04913_ vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__a221o_1
Xhold1333 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2747 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1344 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2758 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1355 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net2769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1366 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1377 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2791 sky130_fd_sc_hd__dlygate4sd3_1
X_08777_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[19\]
+ net656 net602 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout742_A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1388 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 net2802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1399 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2813 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12644__A0 _03623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11447__A1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10655__C1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08863__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13612__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout628_X net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10670_ _05509_ _05950_ vssd1 vssd1 vccd1 vccd1 _06673_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09329_ _05375_ vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_11_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08615__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09748__D net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12340_ _08015_ net355 _03633_ _03634_ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_170_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12271_ _03565_ _03555_ _07951_ vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_33_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14010_ _03879_ _03880_ _03858_ vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_79_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11222_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[37\] _07120_
+ _07184_ _07185_ vssd1 vssd1 vccd1 vccd1 _07186_ sky130_fd_sc_hd__a211o_1
XANTENNA__13059__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11153_ _07094_ _07112_ vssd1 vssd1 vccd1 vccd1 _07119_ sky130_fd_sc_hd__nor2_4
X_10104_ _06128_ _06131_ net513 vssd1 vssd1 vccd1 vccd1 _06132_ sky130_fd_sc_hd__mux2_1
X_11084_ _07043_ _07047_ _07048_ _07050_ vssd1 vssd1 vccd1 vccd1 _07051_ sky130_fd_sc_hd__a31o_1
X_15961_ net1271 vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__inv_2
XANTENNA__12898__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1082 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17700_ clknet_leaf_93_wb_clk_i _03043_ _01396_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[74\]
+ sky130_fd_sc_hd__dfrtp_1
X_10035_ net369 net348 vssd1 vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__nor2_1
X_14912_ net1195 vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__inv_2
X_15892_ net1299 vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_125_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17631_ clknet_leaf_46_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.next_state\[2\]
+ _01327_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14843_ net1176 vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17562_ clknet_leaf_49_wb_clk_i net558 _01258_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write
+ sky130_fd_sc_hd__dfrtp_1
X_14774_ net1101 vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__inv_2
X_11986_ _07796_ _07780_ _07542_ net356 vssd1 vssd1 vccd1 vccd1 _07798_ sky130_fd_sc_hd__o2bb2a_4
XANTENNA__09500__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16513_ clknet_leaf_148_wb_clk_i _02143_ _00209_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13725_ net901 _06918_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[25\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_156_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10937_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[24\] net565 _06925_
+ _06926_ vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__a22o_1
X_17493_ clknet_leaf_38_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[28\]
+ _01189_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08854__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[18\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12927__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13522__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16444_ clknet_leaf_156_wb_clk_i _02074_ _00140_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13656_ net2545 net327 net389 vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__mux2_1
X_10868_ _06808_ _06864_ vssd1 vssd1 vccd1 vccd1 _06865_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17498__Q team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_72_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_116_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12607_ _03650_ net1913 net203 vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__mux2_1
X_16375_ clknet_leaf_146_wb_clk_i _02005_ _00071_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13587_ net2723 net329 net398 vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08606__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10799_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[21\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[21\]
+ vssd1 vssd1 vccd1 vccd1 _06796_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18114_ clknet_leaf_55_wb_clk_i _03437_ _01810_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[31\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_82_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15326_ net1063 vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12538_ net1647 _03650_ net208 vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11610__B2 _07475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18045_ net1037 _03383_ _01741_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.data_from_keypad\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13758__A _05212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15257_ net1057 vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__inv_2
X_12469_ net1765 _03650_ net213 vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__mux2_1
X_14208_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[10\] _04008_
+ net728 vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__a21boi_1
X_15188_ net1069 vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__inv_2
XANTENNA__09674__C net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08204__X _04287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09031__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14139_ net1791 net502 net911 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[22\]
+ sky130_fd_sc_hd__and3_1
Xfanout409 _03728_ vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08700_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[22\]
+ net622 net596 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[22\]
+ _04760_ vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_33_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12601__S _03680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09680_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[1\]
+ net883 net871 net867 vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__and4_1
Xclkbuf_leaf_143_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_143_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08631_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[24\]
+ net838 _04704_ _04705_ vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_85_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17829_ clknet_leaf_103_wb_clk_i _03172_ _01525_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11725__B _07447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12626__A0 _03614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08562_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[25\]
+ net692 net681 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__a22o_1
XANTENNA__09098__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10637__C1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12396__X _03666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08493_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[27\]
+ net645 net615 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[27\]
+ _04556_ vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__a221o_1
XANTENNA__08845__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13432__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout323_A _06737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1065_A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09568__D _04418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09114_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[12\]
+ net818 net806 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__a22o_1
XANTENNA__11601__A1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11601__B2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[23\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09270__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09045_ _05102_ _05103_ vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__nor2_4
XANTENNA_fanout1232_A net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16044__A net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout209_X net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold430 net163 vssd1 vssd1 vccd1 vccd1 net1844 sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[64\] vssd1 vssd1
+ vccd1 vccd1 net1855 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09022__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold452 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[125\] vssd1 vssd1
+ vccd1 vccd1 net1866 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout692_A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold463 net147 vssd1 vssd1 vccd1 vccd1 net1877 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold474 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[76\] vssd1 vssd1
+ vccd1 vccd1 net1888 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10092__A net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold485 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[123\] vssd1 vssd1
+ vccd1 vccd1 net1899 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1020_X net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold496 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[7\] vssd1
+ vssd1 vccd1 vccd1 net1910 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_117_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout910 _03798_ vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__clkbuf_4
Xfanout921 _05213_ vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09881__A _04573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09947_ _05883_ _05975_ vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__or2_1
Xfanout932 net934 vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__buf_2
XANTENNA_fanout480_X net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout943 _04364_ vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__clkbuf_2
Xfanout954 net955 vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout957_A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_146_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout965 net966 vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__buf_4
XANTENNA__13607__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12511__S net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout976 net977 vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__clkbuf_2
Xfanout987 net988 vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__buf_2
X_09878_ _04678_ _05906_ _04637_ vssd1 vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__o21a_1
Xfanout998 net999 vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_5_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1130 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2544 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1141 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net2555 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11635__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08829_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[18\]
+ net664 _04897_ net719 vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__a211o_1
Xhold1152 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2566 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1163 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2577 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1174 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2588 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout745_X net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10340__B2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1185 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 net2599 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1196 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2610 sky130_fd_sc_hd__dlygate4sd3_1
X_11840_ _07651_ _07625_ _07621_ vssd1 vssd1 vccd1 vccd1 _07652_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_16_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13850__B net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08297__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout912_X net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11771_ _07565_ _07572_ vssd1 vssd1 vccd1 vccd1 _07583_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_120_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08836__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13342__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13510_ net2199 net270 net404 vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10722_ _05668_ _06721_ net511 _05669_ vssd1 vssd1 vccd1 vccd1 _06722_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_27_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14490_ net1062 vssd1 vssd1 vccd1 vccd1 _00120_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_172_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13441_ net2137 net264 net413 vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__mux2_1
X_10653_ _05953_ _06656_ net890 vssd1 vssd1 vccd1 vccd1 _06657_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16160_ net1165 vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13372_ net2218 net248 net421 vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__mux2_1
X_10584_ net889 _06591_ net556 vssd1 vssd1 vccd1 vccd1 _06592_ sky130_fd_sc_hd__a21o_1
Xclkload19 clknet_leaf_204_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload19/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__09261__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_156_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_35_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15111_ net1104 vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12323_ _07477_ _03617_ _08022_ _07870_ vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__a211o_1
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16091_ net1308 vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_118_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09775__B _05596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09549__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15042_ net1217 vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__inv_2
X_12254_ _03544_ _03548_ _03512_ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09013__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13896__A2 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11205_ _07086_ _07114_ _07168_ vssd1 vssd1 vccd1 vccd1 _07169_ sky130_fd_sc_hd__and3_2
X_12185_ _07936_ _07940_ _07996_ vssd1 vssd1 vccd1 vccd1 _07997_ sky130_fd_sc_hd__a21oi_2
X_11136_ _07068_ _07071_ _07073_ vssd1 vssd1 vccd1 vccd1 _07102_ sky130_fd_sc_hd__and3_4
XPHY_EDGE_ROW_79_Left_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16993_ clknet_leaf_149_wb_clk_i _02623_ _00689_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13517__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11067_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[1\] team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[0\]
+ vssd1 vssd1 vccd1 vccd1 _07034_ sky130_fd_sc_hd__or2_1
XANTENNA__12421__S net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15944_ net1265 vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__inv_2
XANTENNA__11545__B _07404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10018_ _06040_ _06046_ net530 vssd1 vssd1 vccd1 vccd1 _06047_ sky130_fd_sc_hd__mux2_1
X_15875_ net1304 vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17614_ clknet_leaf_49_wb_clk_i _02985_ _01310_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14826_ net1122 vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__inv_2
XANTENNA__13760__B _06219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17545_ clknet_leaf_49_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[16\]
+ _01241_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14757_ net1184 vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__inv_2
XANTENNA__13281__A0 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11969_ _07741_ _07744_ vssd1 vssd1 vccd1 vccd1 _07781_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12657__A team_05_WB.instance_to_wrap.total_design.core.instr_fetch vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10729__X _06729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13252__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13708_ net901 _06623_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[8\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_195_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_88_Left_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17476_ clknet_leaf_40_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[11\]
+ _01172_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_14688_ net1196 vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16427_ clknet_leaf_185_wb_clk_i _02057_ _00123_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13639_ net2660 net265 net388 vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16358_ clknet_leaf_117_wb_clk_i _01988_ _00054_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10398__A1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15309_ net1082 vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16289_ net1254 vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__inv_2
XANTENNA__09685__B net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08460__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11500__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_11__f_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18028_ clknet_leaf_97_wb_clk_i _03367_ _01724_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire379_X net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09004__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13775__X _03748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_97_Left_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout206 net207 vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__clkbuf_2
Xfanout217 _03660_ vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__buf_4
X_09801_ _05123_ _05144_ vssd1 vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout228 net229 vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_157_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout239 net241 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_52_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09732_ _05760_ _05761_ net585 net583 vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__and4_1
XFILLER_0_66_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08515__A1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09206__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[22\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09663_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[1\]
+ net790 net741 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__a22oi_1
XANTENNA_fanout273_A _06518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08614_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[24\]
+ net673 net666 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09594_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[2\]
+ net786 _05601_ _05610_ _05622_ vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_89_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08545_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[26\]
+ net852 net797 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[26\]
+ _04621_ vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__a221o_1
XFILLER_0_166_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout440_A _03716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14365__B1_N _04092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1182_A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08818__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13162__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08476_ _04533_ _04553_ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__nand2_2
XFILLER_0_77_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09579__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09491__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout705_A _04292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_40_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09243__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08451__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12506__S net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09028_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[14\]
+ net797 net780 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout695_X net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold260 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[6\] vssd1 vssd1
+ vccd1 vccd1 net1674 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[4\] vssd1 vssd1
+ vccd1 vccd1 net1685 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold282 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[119\] vssd1 vssd1
+ vccd1 vccd1 net1696 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold293 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[24\] vssd1 vssd1
+ vccd1 vccd1 net1707 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout862_X net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout740 _04421_ vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13337__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout751 _04415_ vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__buf_4
XANTENNA__15118__A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout762 net763 vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__buf_4
X_13990_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[6\] _03840_ _03843_
+ vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__a21oi_1
Xfanout773 _04406_ vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__buf_4
Xfanout784 net785 vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__buf_4
Xfanout795 _04395_ vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__buf_4
X_12941_ net252 net2852 net468 vssd1 vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_161_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15660_ net1282 vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__inv_2
X_12872_ net247 net2273 net477 vssd1 vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__mux2_1
X_14611_ net1216 vssd1 vssd1 vccd1 vccd1 _00241_ sky130_fd_sc_hd__inv_2
X_11823_ _07633_ _07634_ _07619_ vssd1 vssd1 vccd1 vccd1 _07635_ sky130_fd_sc_hd__a21oi_2
X_15591_ net1249 vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__inv_2
XANTENNA__08809__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[19\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13072__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10077__B1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17330_ clknet_leaf_125_wb_clk_i _02960_ _01026_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_14542_ net1184 vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__inv_2
X_11754_ _07553_ _07558_ vssd1 vssd1 vccd1 vccd1 _07566_ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09482__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_7__f_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15788__A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17261_ clknet_leaf_161_wb_clk_i _02891_ _00957_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10705_ _05804_ _05806_ vssd1 vssd1 vccd1 vccd1 _06706_ sky130_fd_sc_hd__xnor2_4
X_14473_ net1222 vssd1 vssd1 vccd1 vccd1 _00103_ sky130_fd_sc_hd__inv_2
X_11685_ net52 net51 net54 net53 vssd1 vssd1 vccd1 vccd1 _07499_ sky130_fd_sc_hd__or4_1
XANTENNA__08690__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16212_ net1061 vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09786__A net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13424_ net2876 net321 net416 vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__mux2_1
X_10636_ _05423_ _05814_ vssd1 vssd1 vccd1 vccd1 _06641_ sky130_fd_sc_hd__xor2_2
XFILLER_0_24_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17192_ clknet_leaf_203_wb_clk_i _02822_ _00888_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload108 clknet_leaf_160_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload108/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16143_ net1273 vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload119 clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload119/Y sky130_fd_sc_hd__inv_6
XFILLER_0_23_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08442__B1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13355_ net316 net2838 net427 vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__mux2_1
XANTENNA__12416__S net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10567_ net889 _06572_ _06575_ net554 vssd1 vssd1 vccd1 vccd1 _06576_ sky130_fd_sc_hd__a211o_1
XFILLER_0_12_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12306_ _03596_ _03598_ _03599_ _03600_ vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__or4_2
X_16074_ net1174 vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13286_ net295 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[8\]
+ net435 vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__mux2_1
X_10498_ _05058_ _05923_ _06507_ _06510_ _06060_ vssd1 vssd1 vccd1 vccd1 _06511_ sky130_fd_sc_hd__o32a_1
X_15025_ net1192 vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__inv_2
X_12237_ _08015_ _03529_ vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13755__B _06350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12168_ _07932_ _07968_ _07977_ vssd1 vssd1 vccd1 vccd1 _07980_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11556__A _07379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13247__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11119_ _07082_ _07084_ _07085_ vssd1 vssd1 vccd1 vccd1 _07086_ sky130_fd_sc_hd__nor3_1
XANTENNA__12004__X _07816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16976_ clknet_leaf_138_wb_clk_i _02606_ _00672_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_12099_ _07902_ _07910_ vssd1 vssd1 vccd1 vccd1 _07911_ sky130_fd_sc_hd__and2_1
XANTENNA__09671__D net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput6 DAT_I[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
X_15927_ net1294 vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_3_4_0_wb_clk_i_X clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15858_ net1299 vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14809_ net1053 vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__inv_2
X_15789_ net1270 vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08330_ net948 net937 net933 vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17528_ clknet_leaf_109_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[31\]
+ _01224_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[31\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10607__A2 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09473__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08261_ net968 net953 _04269_ vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__or3_4
XFILLER_0_74_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11280__A2 _07105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17459_ clknet_leaf_66_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[27\]
+ _01155_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_144_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08192_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[13\] _04274_
+ _04239_ vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__a21oi_4
XANTENNA__09225__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10635__A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08599__X team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[25\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout390_A _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13157__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout488_A _03700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11466__A _07352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10370__A net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09581__D net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09715_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[0\]
+ net951 net931 net926 vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__and4_1
XANTENNA__12996__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09646_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[1\]
+ net940 net1013 net927 vssd1 vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__and4_1
XFILLER_0_69_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09577_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[2\]
+ net947 net935 net924 vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout822_A net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout443_X net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08528_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[26\]
+ net619 net596 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09464__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[5\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11271__A2 _07103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08672__B1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout610_X net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08459_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[28\]
+ net803 net740 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout708_X net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13620__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15401__A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11470_ net1050 net1049 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[0\]
+ vssd1 vssd1 vccd1 vccd1 _07381_ sky130_fd_sc_hd__o21a_1
XFILLER_0_135_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09216__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10421_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[18\] _06095_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[19\]
+ vssd1 vssd1 vccd1 vccd1 _06438_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08424__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13140_ net256 net2789 net445 vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__mux2_1
X_10352_ net1020 _04798_ _04799_ vssd1 vssd1 vccd1 vccd1 _06372_ sky130_fd_sc_hd__o21ai_1
X_13071_ net228 net2552 net453 vssd1 vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__mux2_1
X_10283_ _06075_ _06077_ vssd1 vssd1 vccd1 vccd1 _06306_ sky130_fd_sc_hd__nor2_1
X_12022_ _07773_ _07775_ _07815_ _07833_ vssd1 vssd1 vccd1 vccd1 _07834_ sky130_fd_sc_hd__o31a_1
XANTENNA_input49_A wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_163_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_10__f_wb_clk_i_X clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13067__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16830_ clknet_leaf_163_wb_clk_i _02460_ _00526_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout570 _04344_ vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__buf_4
Xfanout581 net582 vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__clkbuf_2
Xfanout592 _04368_ vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__buf_6
X_13973_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[10\] _03844_ vssd1
+ vssd1 vccd1 vccd1 _03845_ sky130_fd_sc_hd__and2_1
X_16761_ clknet_leaf_9_wb_clk_i _02391_ _00457_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_15712_ net1153 vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__inv_2
X_12924_ net323 net1876 net472 vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__mux2_1
X_16692_ clknet_leaf_112_wb_clk_i _02322_ _00388_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12855_ net313 net2259 net482 vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__mux2_1
X_15643_ net1245 vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__inv_2
X_11806_ _07610_ _07611_ _07617_ vssd1 vssd1 vccd1 vccd1 _07618_ sky130_fd_sc_hd__a21oi_1
X_18362_ net1347 vssd1 vssd1 vccd1 vccd1 la_data_out[10] sky130_fd_sc_hd__buf_2
XFILLER_0_68_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15574_ net1247 vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12786_ net320 net2355 net488 vssd1 vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09455__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17313_ clknet_leaf_150_wb_clk_i _02943_ _01009_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[9\]
+ sky130_fd_sc_hd__dfrtp_2
X_14525_ net1089 vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__inv_2
XANTENNA__11262__A2 _07091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11737_ _07534_ _07539_ _07543_ _07544_ vssd1 vssd1 vccd1 vccd1 _07549_ sky130_fd_sc_hd__o22a_1
XFILLER_0_56_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18293_ net1385 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
XANTENNA__08663__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13530__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17244_ clknet_leaf_156_wb_clk_i _02874_ _00940_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14456_ net1207 vssd1 vssd1 vccd1 vccd1 _00086_ sky130_fd_sc_hd__inv_2
X_11668_ net13 net991 net918 net2731 vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13407_ net2247 net257 net416 vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__mux2_1
XANTENNA__11014__A2 _06768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10619_ net894 _06622_ _06624_ vssd1 vssd1 vccd1 vccd1 _06625_ sky130_fd_sc_hd__a21o_1
X_17175_ clknet_leaf_147_wb_clk_i _02805_ _00871_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08415__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14387_ net1550 vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11599_ net1618 net1009 net346 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16126_ net1136 vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13338_ net228 net2786 net426 vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16057_ net1262 vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__inv_2
X_13269_ net239 net2585 net434 vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15008_ net1102 vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__inv_2
XANTENNA__09682__C net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10190__A _04265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18344__1333 vssd1 vssd1 vccd1 vccd1 _18344__1333/HI net1333 sky130_fd_sc_hd__conb_1
XFILLER_0_138_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13475__A0 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16959_ clknet_leaf_153_wb_clk_i _02589_ _00655_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_09500_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[4\]
+ net649 net603 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[4\]
+ _05534_ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__a221o_1
XANTENNA__10289__B1 _04275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09694__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09431_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[5\]
+ net678 net635 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[5\]
+ _05473_ vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__a221o_1
XANTENNA__13227__A0 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18359__1344 vssd1 vssd1 vccd1 vccd1 _18359__1344/HI net1344 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09362_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[7\]
+ net796 net739 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05408_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_47_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09446__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08313_ net950 net936 net929 vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__and3_2
XFILLER_0_157_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12450__A1 _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08654__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09293_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[8\]
+ net714 net654 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__a22o_1
XANTENNA_11 _07410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13440__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout236_A net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08244_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[31\]
+ net630 net599 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_43_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11005__A2 _06572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08175_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[11\] _04249_
+ vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__nand2_2
XANTENNA_clkbuf_4_6__f_wb_clk_i_X clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10365__A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09576__D net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput140 net140 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1312_A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput151 net151 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput162 net162 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
Xoutput173 net173 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__clkbuf_4
Xoutput184 net184 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout772_A _04406_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout393_X net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11483__X _07394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout658_X net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11924__A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13615__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10970_ _06804_ _06805_ _06867_ vssd1 vssd1 vccd1 vccd1 _06953_ sky130_fd_sc_hd__o21ai_1
XANTENNA__14300__A net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09629_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[2\]
+ net633 _05663_ net720 vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_67_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08893__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout825_X net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12640_ net1776 _07816_ _03682_ vssd1 vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_139_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09437__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12571_ net1754 _07821_ _03678_ vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__mux2_1
XANTENNA__12441__A1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08645__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13350__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14310_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[16\] _04990_
+ _04965_ _04944_ vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_156_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11522_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[15\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[15\]
+ net1031 vssd1 vssd1 vccd1 vccd1 _07433_ sky130_fd_sc_hd__mux2_1
XANTENNA__15131__A net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15290_ net1062 vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14241_ team_05_WB.instance_to_wrap.total_design.keypad0.counter\[7\] _04020_ net2524
+ vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__a21oi_1
X_11453_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[3\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[3\]
+ net1035 vssd1 vssd1 vccd1 vccd1 _07364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08948__A1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10404_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[20\] net903 _06418_
+ _06421_ vssd1 vssd1 vccd1 vccd1 _06422_ sky130_fd_sc_hd__a211o_2
XFILLER_0_21_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14172_ net1942 net506 net909 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[21\]
+ sky130_fd_sc_hd__and3_1
X_11384_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[3\] _07314_
+ vssd1 vssd1 vccd1 vccd1 _07315_ sky130_fd_sc_hd__nand2_1
XANTENNA__09070__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13123_ net309 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[3\]
+ net448 vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__mux2_1
X_10335_ _05929_ net510 _06355_ _06017_ _06354_ vssd1 vssd1 vccd1 vccd1 _06356_ sky130_fd_sc_hd__o221a_1
X_17931_ clknet_leaf_43_wb_clk_i _03270_ _01627_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13054_ net317 net2371 net457 vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__mux2_1
X_10266_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[26\] _06100_ vssd1
+ vssd1 vccd1 vccd1 _06290_ sky130_fd_sc_hd__nor2_1
Xfanout1310 net1311 vssd1 vssd1 vccd1 vccd1 net1310 sky130_fd_sc_hd__buf_2
X_12005_ _07773_ _07776_ vssd1 vssd1 vccd1 vccd1 _07817_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17862_ clknet_leaf_76_wb_clk_i _03205_ _01558_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10197_ _06115_ _06123_ net517 vssd1 vssd1 vccd1 vccd1 _06223_ sky130_fd_sc_hd__mux2_1
X_16813_ clknet_leaf_162_wb_clk_i _02443_ _00509_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_17793_ clknet_leaf_100_wb_clk_i _03136_ _01489_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[103\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13525__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16744_ clknet_leaf_1_wb_clk_i _02374_ _00440_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13956_ _03826_ _03827_ vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09304__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[20\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12907_ net255 net2172 net472 vssd1 vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__mux2_1
X_13887_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[15\]
+ net560 net576 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[15\]
+ net987 vssd1 vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__a221o_1
X_16675_ clknet_leaf_192_wb_clk_i _02305_ _00371_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08884__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15626_ net1159 vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__inv_2
X_12838_ net227 net2621 net481 vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09428__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18345_ net34 vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12432__A1 _07821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11235__A2 _07113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15557_ net1118 vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__inv_2
X_12769_ net232 net2924 net490 vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__mux2_1
XANTENNA__08636__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08100__A2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[11\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13260__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_168_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_168_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_14508_ net1109 vssd1 vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__inv_2
X_15488_ net1154 vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__inv_2
X_18276_ clknet_leaf_36_wb_clk_i _03505_ _01971_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_126_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09677__C net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10994__A1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput20 DAT_I[26] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
X_17227_ clknet_leaf_160_wb_clk_i _02857_ _00923_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput31 DAT_I[7] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14439_ net1105 vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput42 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput53 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_1
Xinput64 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold804 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2218 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09061__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17158_ clknet_leaf_119_wb_clk_i _02788_ _00854_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold815 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2229 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10746__A1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold826 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold837 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2251 sky130_fd_sc_hd__dlygate4sd3_1
X_16109_ net1152 vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__inv_2
Xhold848 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2262 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12604__S net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17089_ clknet_leaf_148_wb_clk_i _02719_ _00785_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09980_ _06005_ _06008_ net516 vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold859 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2273 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08931_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[16\]
+ net833 net826 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__a22o_1
XANTENNA__12499__A1 _03605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10632__B _06637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08862_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[17\]
+ net700 net602 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__a22o_1
Xhold1504 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2918 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08877__X _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1515 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net2929 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1526 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2940 sky130_fd_sc_hd__dlygate4sd3_1
X_08793_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[19\]
+ net810 net737 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__a22o_1
Xhold1537 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net2951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1548 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net2962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1559 team_05_WB.instance_to_wrap.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 net2973
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13435__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09667__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11474__A2 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08875__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout353_A _03717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09414_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[6\]
+ net838 net757 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_45_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09419__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09345_ _05385_ _05387_ _05389_ _05391_ vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__or4_1
XFILLER_0_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12423__A1 _07812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11226__A2 _07099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08627__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout520_A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16047__A net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout618_A net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13170__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Left_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09276_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[9\]
+ net776 net734 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_134_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08227_ net884 net872 net858 vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1050_X net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout406_X net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08158_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[4\] team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__nand2b_4
XANTENNA__09052__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout987_A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12514__S _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08089_ net1023 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__and2b_1
X_10120_ _06144_ _06147_ net513 vssd1 vssd1 vccd1 vccd1 _06148_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout775_X net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_42_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10051_ _06076_ _06079_ net514 vssd1 vssd1 vccd1 vccd1 _06080_ sky130_fd_sc_hd__mux2_1
XANTENNA__13853__B net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13345__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13810_ net1597 net969 net724 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[21\]
+ sky130_fd_sc_hd__and3_1
X_14790_ net1208 vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13741_ net923 _06609_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[9\]
+ sky130_fd_sc_hd__nor2_1
X_10953_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[21\] net567 _06938_
+ _06939_ vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_27_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08866__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16460_ clknet_leaf_7_wb_clk_i _02090_ _00156_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13672_ net2424 net265 net384 vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__mux2_1
X_10884_ _06784_ _06880_ vssd1 vssd1 vccd1 vccd1 _06881_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_51_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12623_ _03610_ net1873 net202 vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__mux2_1
X_15411_ net1133 vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_62_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11217__A2 _07100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16391_ clknet_leaf_203_wb_clk_i _02021_ _00087_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13080__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18130_ clknet_leaf_48_wb_clk_i _00026_ _01826_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10425__B1 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15342_ net1187 vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__inv_2
X_12554_ _03655_ net1796 net206 vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09291__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18343__1332 vssd1 vssd1 vccd1 vccd1 _18343__1332/HI net1332 sky130_fd_sc_hd__conb_1
XFILLER_0_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10717__B team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09830__A2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11505_ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[10\] _07415_ net1002
+ vssd1 vssd1 vccd1 vccd1 _07416_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15796__A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18061_ clknet_leaf_98_wb_clk_i _03399_ _01757_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__dfrtp_1
X_15273_ net1221 vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12485_ net1794 _03655_ net210 vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14224_ team_05_WB.instance_to_wrap.total_design.keypad0.counter\[6\] _04019_ vssd1
+ vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__and2_1
XANTENNA__09794__A _05208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17012_ clknet_leaf_120_wb_clk_i _02642_ _00708_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11436_ team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.state\[1\] team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.state\[2\]
+ team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.state\[0\] vssd1 vssd1 vccd1
+ vccd1 _07349_ sky130_fd_sc_hd__or3b_4
XFILLER_0_111_418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08397__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14155_ _03859_ net907 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[4\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12424__S _03667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11367_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[0\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[0\]
+ _06839_ _06840_ vssd1 vssd1 vccd1 vccd1 _07306_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18358__1343 vssd1 vssd1 vccd1 vccd1 _18358__1343/HI net1343 sky130_fd_sc_hd__conb_1
X_13106_ net252 net2873 net448 vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_60_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10318_ _06003_ _06329_ _06332_ _06339_ vssd1 vssd1 vccd1 vccd1 _06340_ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14086_ _03932_ _03952_ vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__nor2_1
X_11298_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[65\] _07118_
+ _07256_ _07257_ vssd1 vssd1 vccd1 vccd1 _07258_ sky130_fd_sc_hd__a211o_1
X_17914_ clknet_leaf_63_wb_clk_i _03257_ _01610_ vssd1 vssd1 vccd1 vccd1 team_05_WB.EN_VAL_REG
+ sky130_fd_sc_hd__dfrtp_4
X_13037_ net233 net2461 net459 vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__mux2_1
X_10249_ _05907_ _06272_ vssd1 vssd1 vccd1 vccd1 _06273_ sky130_fd_sc_hd__and2b_2
XFILLER_0_28_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1140 net1141 vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__buf_4
Xfanout1151 net1177 vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__clkbuf_2
Xfanout1162 net1163 vssd1 vssd1 vccd1 vccd1 net1162 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13763__B _05921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17845_ clknet_leaf_91_wb_clk_i _03188_ _01541_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[91\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1173 net1174 vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__buf_4
Xfanout1184 net1186 vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__buf_4
XANTENNA__13255__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1195 net1198 vssd1 vssd1 vccd1 vccd1 net1195 sky130_fd_sc_hd__buf_4
X_17776_ clknet_leaf_93_wb_clk_i _03119_ _01472_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14988_ net1111 vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16727_ clknet_leaf_150_wb_clk_i _02357_ _00423_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13939_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[5\] team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14875__A net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10664__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16658_ clknet_leaf_125_wb_clk_i _02288_ _00354_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15609_ net1168 vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__inv_2
XANTENNA__11208__A2 _07103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08609__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16589_ clknet_leaf_160_wb_clk_i _02219_ _00285_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11503__S net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09130_ net572 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[12\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[12\] vssd1 vssd1 vccd1
+ vccd1 _05185_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_174_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18328_ team_05_WB.instance_to_wrap.lcd_rs vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09821__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09061_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[13\]
+ net712 net683 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[13\]
+ _05105_ vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18259_ clknet_leaf_40_wb_clk_i _03488_ _01954_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_170_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09034__B1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold601 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2015 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10914__Y _06907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold612 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2026 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold623 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 net2037 sky130_fd_sc_hd__dlygate4sd3_1
Xhold634 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2048 sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2059 sky130_fd_sc_hd__dlygate4sd3_1
Xhold656 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2070 sky130_fd_sc_hd__dlygate4sd3_1
Xhold667 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 net2081 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_107_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09963_ _04636_ _05902_ _05990_ _05928_ vssd1 vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold678 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net2092 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold689 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net2103 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_65_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08914_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[16\]
+ net703 net695 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[16\]
+ _04978_ vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1010_A net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09894_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[14\] _04272_
+ vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__nand2_4
XANTENNA_fanout1108_A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1301 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 net2715 sky130_fd_sc_hd__dlygate4sd3_1
X_08845_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[18\]
+ net818 net790 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__a22o_1
Xhold1312 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2726 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1323 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net2737 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout470_A net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1334 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2748 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1345 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2759 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13165__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout568_A _06774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1356 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 net2770 sky130_fd_sc_hd__dlygate4sd3_1
X_08776_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[19\]
+ net652 net594 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[19\]
+ _04842_ vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__a221o_1
Xhold1367 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1378 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net2792 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1389 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net2803 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_108_Left_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11447__A2 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08848__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout735_A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout902_A _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09328_ _05351_ _05374_ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_153_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09273__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09812__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09259_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[21\] net967
+ _04246_ _04352_ vssd1 vssd1 vccd1 vccd1 _05310_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_clkbuf_leaf_146_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_8_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_170_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_117_Left_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12270_ _07969_ _03556_ vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09025__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout892_X net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11221_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[37\] _07097_
+ _07119_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[29\] _07031_
+ vssd1 vssd1 vccd1 vccd1 _07185_ sky130_fd_sc_hd__a221o_1
XANTENNA__08379__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12580__A0 _03661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11152_ _07074_ _07114_ vssd1 vssd1 vccd1 vccd1 _07118_ sky130_fd_sc_hd__nor2_4
X_10103_ _06129_ _06130_ vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__nand2_1
X_11083_ _07046_ _07049_ vssd1 vssd1 vccd1 vccd1 _07050_ sky130_fd_sc_hd__nand2_1
X_15960_ net1266 vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input31_A DAT_I[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10034_ _05531_ _06061_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__or2_1
X_14911_ net1179 vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15891_ net1303 vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__inv_2
XANTENNA__13075__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17630_ clknet_leaf_51_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.next_state\[1\]
+ _01326_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08551__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14842_ net1053 vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_125_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17561_ clknet_leaf_49_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.next_read
+ _01257_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__12635__A1 _07797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11985_ _07796_ _07782_ _07553_ net356 vssd1 vssd1 vccd1 vccd1 _07797_ sky130_fd_sc_hd__o2bb2a_4
X_14773_ net1060 vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__inv_2
XANTENNA__08839__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08303__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10646__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16512_ clknet_leaf_127_wb_clk_i _02142_ _00208_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13724_ net900 _06320_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[24\]
+ sky130_fd_sc_hd__nor2_1
X_10936_ net960 _06320_ net565 vssd1 vssd1 vccd1 vccd1 _06926_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_169_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17492_ clknet_leaf_36_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[27\]
+ _01188_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_185_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_156_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16443_ clknet_leaf_189_wb_clk_i _02073_ _00139_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12419__S net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10867_ _06812_ _06862_ _06810_ vssd1 vssd1 vccd1 vccd1 _06864_ sky130_fd_sc_hd__a21oi_2
X_13655_ net2115 net322 net389 vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12606_ net1741 _07816_ _03680_ vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16374_ clknet_leaf_150_wb_clk_i _02004_ _00070_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09264__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13586_ net2942 net316 net399 vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__mux2_1
X_10798_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[21\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[21\]
+ vssd1 vssd1 vccd1 vccd1 _06795_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18113_ clknet_leaf_69_wb_clk_i _03436_ _01809_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[30\]
+ sky130_fd_sc_hd__dfrtp_2
X_12537_ _07816_ net1809 _03675_ vssd1 vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__mux2_1
XANTENNA__12365__D _03659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15325_ net1090 vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11610__A2 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18044_ clknet_leaf_54_wb_clk_i _03382_ _01740_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_12468_ net1970 _07816_ _03670_ vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__mux2_1
XANTENNA__13758__B _06273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15256_ net1243 vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12662__B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14207_ _04008_ net728 _04007_ vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__and3b_1
X_11419_ net1926 _07323_ vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__xor2_1
XFILLER_0_151_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15187_ net1213 vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__inv_2
X_12399_ net1685 _07816_ _07852_ vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__mux2_1
XANTENNA__09674__D net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14138_ net1942 net506 net911 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[21\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_10_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08790__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14069_ _03936_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[11\] _03935_
+ vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08630_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[24\]
+ net783 net761 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__a22o_1
XANTENNA__08542__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17828_ clknet_leaf_80_wb_clk_i _03171_ _01524_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_146_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11725__C _07478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08561_ _04636_ vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17759_ clknet_leaf_88_wb_clk_i _03102_ _01455_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_183_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_183_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_18_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09699__A _05731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08492_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[27\]
+ net708 _04569_ net721 vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__a211o_1
XFILLER_0_49_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_112_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_112_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09113_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[12\]
+ net814 net802 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[12\]
+ _05168_ vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11601__A2 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1058_A net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09044_ _05078_ _05100_ vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09007__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold420 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[88\] vssd1 vssd1
+ vccd1 vccd1 net1834 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold431 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[27\] vssd1 vssd1
+ vccd1 vccd1 net1845 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09584__D net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold442 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[49\] vssd1 vssd1
+ vccd1 vccd1 net1856 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1225_A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold453 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[102\] vssd1 vssd1
+ vccd1 vccd1 net1867 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1034 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold464 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[119\] vssd1 vssd1
+ vccd1 vccd1 net1878 sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[47\] vssd1 vssd1
+ vccd1 vccd1 net1889 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12999__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold486 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[1\] vssd1 vssd1
+ vccd1 vccd1 net1900 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout900 net902 vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout685_A net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold497 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[40\] vssd1 vssd1
+ vccd1 vccd1 net1911 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout911 net912 vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout922 _05213_ vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08781__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09946_ _05930_ _05974_ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_74_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout933 net934 vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1013_X net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout944 _04364_ vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__buf_2
Xfanout955 _04245_ vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__buf_2
Xfanout966 net967 vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_146_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout977 _04178_ vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11668__A2 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ _04717_ _05899_ _05904_ vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__a21oi_1
Xhold1120 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net2534 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout473_X net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout852_A _04370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout988 _03762_ vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__buf_2
X_18342__1331 vssd1 vssd1 vccd1 vccd1 _18342__1331/HI net1331 sky130_fd_sc_hd__conb_1
Xfanout999 net1000 vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1131 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net2545 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08533__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1142 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2556 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08828_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[18\]
+ net640 net598 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__a22o_1
Xhold1153 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1164 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2578 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1175 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net2589 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1186 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net2600 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12617__A1 _07789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08759_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[21\]
+ net803 net746 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__a22o_1
Xhold1197 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2611 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout640_X net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout738_X net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13623__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10628__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11770_ _07569_ _07581_ vssd1 vssd1 vccd1 vccd1 _07582_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_120_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09494__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18357__1342 vssd1 vssd1 vccd1 vccd1 _18357__1342/HI net1342 sky130_fd_sc_hd__conb_1
X_10721_ net1018 _05667_ net551 vssd1 vssd1 vccd1 vccd1 _06721_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_172_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout905_X net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13440_ net2450 net258 net412 vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__mux2_1
X_10652_ _05812_ _05952_ vssd1 vssd1 vccd1 vccd1 _06656_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09246__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_125_Left_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13371_ net2843 net227 net421 vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__mux2_1
X_10583_ _05284_ _05821_ vssd1 vssd1 vccd1 vccd1 _06591_ sky130_fd_sc_hd__xnor2_2
X_12322_ _03616_ vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15110_ net1209 vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16090_ net1308 vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08305__X _04387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15041_ net1236 vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12253_ _08019_ _03543_ vssd1 vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__nand2_1
XANTENNA__12553__A0 _03646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11204_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[4\] _04163_
+ _07061_ _07067_ _07038_ vssd1 vssd1 vccd1 vccd1 _07168_ sky130_fd_sc_hd__a311oi_1
X_12184_ _07931_ _07940_ _07936_ vssd1 vssd1 vccd1 vccd1 _07996_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11135_ _07038_ _07068_ _07079_ vssd1 vssd1 vccd1 vccd1 _07101_ sky130_fd_sc_hd__and3_4
XANTENNA__08772__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12702__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16992_ clknet_leaf_126_wb_clk_i _02622_ _00688_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11066_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[1\] team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[0\]
+ vssd1 vssd1 vccd1 vccd1 _07033_ sky130_fd_sc_hd__nor2_1
X_15943_ net1291 vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__inv_2
XANTENNA__08524__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10017_ _06042_ _06045_ net514 vssd1 vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__mux2_1
X_15874_ net1288 vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__inv_2
X_17613_ clknet_leaf_49_wb_clk_i _02984_ _01309_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12608__A1 _07836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14825_ net1222 vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__inv_2
XANTENNA__13533__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17544_ clknet_leaf_61_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[15\]
+ _01240_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09485__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14756_ net1230 vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__inv_2
X_11968_ _07778_ _07779_ _07529_ vssd1 vssd1 vccd1 vccd1 _07780_ sky130_fd_sc_hd__a21o_1
XFILLER_0_58_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12657__B net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13707_ net900 _06641_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[7\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__11292__B1 _07126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10919_ net961 _06907_ net566 vssd1 vssd1 vccd1 vccd1 _06912_ sky130_fd_sc_hd__a21oi_1
X_17475_ clknet_leaf_41_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[10\]
+ _01171_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14687_ net1178 vssd1 vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11899_ _07672_ _07673_ _07650_ vssd1 vssd1 vccd1 vccd1 _07711_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_920 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16426_ clknet_leaf_196_wb_clk_i _02056_ _00122_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13638_ net2004 net257 net388 vssd1 vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__mux2_1
XANTENNA__09237__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16357_ clknet_leaf_175_wb_clk_i _01987_ _00053_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13569_ net2142 net227 net399 vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12792__A0 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11595__B2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[29\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15308_ net1072 vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16288_ net1254 vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__inv_2
XANTENNA__09685__C net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18027_ clknet_leaf_97_wb_clk_i _03366_ _01723_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_15239_ net1105 vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__inv_2
XFILLER_0_160_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09982__A _05442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17972__Q net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout207 _03679_ vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__clkbuf_4
X_09800_ _05123_ _05144_ vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__nor2_1
XANTENNA__08763__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout218 net221 vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__clkbuf_2
Xfanout229 _06385_ vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_163_Right_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09731_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[0\]
+ net748 _05739_ _05740_ _05742_ vssd1 vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__08515__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[27\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09662_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[1\]
+ _04366_ net815 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[1\]
+ net854 vssd1 vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_94_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08613_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[24\]
+ net623 net616 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[24\]
+ _04687_ vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__a221o_1
X_09593_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[2\]
+ net829 _05611_ _05613_ net853 vssd1 vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_94_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_141_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13443__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08544_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[26\]
+ net848 net735 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__a22o_1
XANTENNA__15224__A net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09476__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08475_ net573 _04552_ _04361_ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10368__A _05886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout433_A _03722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1175_A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09579__D net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout600_A net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout221_X net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_80_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09027_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[14\]
+ net828 net747 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold250 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[6\] vssd1 vssd1
+ vccd1 vccd1 net1664 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold261 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[110\] vssd1 vssd1
+ vccd1 vccd1 net1675 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout590_X net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold272 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[29\]
+ vssd1 vssd1 vccd1 vccd1 net1686 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout688_X net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold283 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[12\] vssd1 vssd1
+ vccd1 vccd1 net1697 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13618__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold294 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[20\] vssd1 vssd1
+ vccd1 vccd1 net1708 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08754__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12522__S net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14303__A _04533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout730 _07320_ vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__clkbuf_2
Xfanout741 net744 vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_165_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09929_ _05285_ _05817_ _05957_ vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__and3_1
Xfanout752 net755 vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08301__A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout763 _04411_ vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__buf_4
Xfanout774 net777 vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__buf_6
XANTENNA_fanout855_X net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08506__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout785 _04401_ vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__buf_4
Xfanout796 net797 vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__clkbuf_8
X_12940_ net246 net2214 net469 vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ net226 net2196 net478 vssd1 vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__mux2_1
XANTENNA__13353__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14610_ net1232 vssd1 vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__inv_2
X_11822_ _07611_ _07630_ vssd1 vssd1 vccd1 vccd1 _07634_ sky130_fd_sc_hd__xnor2_2
X_15590_ net1249 vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__inv_2
XANTENNA__10077__A1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[31\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09132__A _05165_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11274__B1 _07108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10077__B2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[31\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14541_ net1081 vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11753_ net549 _07522_ vssd1 vssd1 vccd1 vccd1 _07565_ sky130_fd_sc_hd__nand2_2
X_10704_ net1969 net330 net540 vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__mux2_1
X_17260_ clknet_leaf_2_wb_clk_i _02890_ _00956_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11684_ _07494_ _07495_ _07496_ _07497_ vssd1 vssd1 vccd1 vccd1 _07498_ sky130_fd_sc_hd__or4_1
X_14472_ net1223 vssd1 vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__inv_2
XANTENNA__09219__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16211_ net1074 vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10635_ net891 _06639_ vssd1 vssd1 vccd1 vccd1 _06640_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13423_ net2452 net311 net416 vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17191_ clknet_leaf_199_wb_clk_i _02821_ _00887_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload109 clknet_leaf_161_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload109/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16142_ net1273 vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13354_ net318 net2548 net424 vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__mux2_1
X_10566_ _06573_ _06574_ net889 vssd1 vssd1 vccd1 vccd1 _06575_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12305_ _03512_ _03583_ vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__nor2_1
XANTENNA__08993__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16073_ net1173 vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__inv_2
X_13285_ net300 net2626 net435 vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__mux2_1
X_10497_ net369 net347 vssd1 vssd1 vccd1 vccd1 _06510_ sky130_fd_sc_hd__or2_2
X_12236_ _03511_ _03524_ _03528_ _03529_ _07992_ vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__a32o_2
XFILLER_0_121_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15024_ net1093 vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13528__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12432__S _03667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12167_ _07968_ _07977_ _07932_ vssd1 vssd1 vccd1 vccd1 _07979_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_9_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11118_ _07052_ _07071_ _07075_ vssd1 vssd1 vccd1 vccd1 _07085_ sky130_fd_sc_hd__and3_1
XANTENNA__11556__B _07465_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16975_ clknet_leaf_134_wb_clk_i _02605_ _00671_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_12098_ _07905_ _07906_ _07907_ _07864_ vssd1 vssd1 vccd1 vccd1 _07910_ sky130_fd_sc_hd__o22ai_4
XTAP_TAPCELL_ROW_30_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15926_ net1257 vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__inv_2
X_11049_ net960 _06706_ net566 vssd1 vssd1 vccd1 vccd1 _07018_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput7 DAT_I[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09170__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15857_ net1270 vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__inv_2
XANTENNA__13263__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14808_ net1244 vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15788_ net1300 vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17527_ clknet_leaf_73_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[30\]
+ _01223_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[30\]
+ sky130_fd_sc_hd__dfrtp_4
X_14739_ net1214 vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08260_ net967 net954 _04269_ vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__nor3_1
XFILLER_0_117_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09977__A _05596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17458_ clknet_leaf_65_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[26\]
+ _01154_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17967__Q net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16409_ clknet_leaf_9_wb_clk_i _02039_ _00105_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08191_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[14\] _04273_
+ vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__nor2_2
XFILLER_0_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17389_ clknet_leaf_58_wb_clk_i net1443 _01085_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12607__S net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11568__A1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11511__S net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18341__1330 vssd1 vssd1 vccd1 vccd1 _18341__1330/HI net1330 sky130_fd_sc_hd__conb_1
XANTENNA__13786__X _03759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08984__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12517__A0 _07793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08736__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13438__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15219__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18356__1341 vssd1 vssd1 vccd1 vccd1 _18356__1341/HI net1341 sky130_fd_sc_hd__conb_1
XFILLER_0_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10370__B _05977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout383_A _04265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09714_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[0\]
+ net951 net936 net934 vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__and4_1
XFILLER_0_97_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09645_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[1\]
+ net946 net932 net930 vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout550_A _07448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13173__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout648_A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09576_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[2\]
+ net940 net935 net927 vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__and4_1
XFILLER_0_96_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09449__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11256__B1 _07129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08527_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[26\]
+ net674 net635 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[26\]
+ _04603_ vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__a221o_1
XFILLER_0_171_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10098__A _05256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout815_A _04388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout436_X net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08458_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[28\]
+ net776 net747 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[28\]
+ _04536_ vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__a221o_1
XFILLER_0_147_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold226_A team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12517__S _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10385__X _06404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08389_ net380 _04466_ vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout603_X net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10420_ _06428_ _06436_ net536 vssd1 vssd1 vccd1 vccd1 _06437_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09621__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10351_ net893 _06368_ _06370_ net555 vssd1 vssd1 vccd1 vccd1 _06371_ sky130_fd_sc_hd__a211o_1
XANTENNA__08975__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13070_ net231 net2407 net454 vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10282_ net524 _06201_ _06304_ vssd1 vssd1 vccd1 vccd1 _06305_ sky130_fd_sc_hd__a21oi_1
X_12021_ _07767_ _07769_ _07773_ _07765_ vssd1 vssd1 vccd1 vccd1 _07833_ sky130_fd_sc_hd__o31ai_1
XANTENNA__13348__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10561__A net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout560 net561 vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__buf_2
XANTENNA__14968__A net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout571 net573 vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__clkbuf_4
Xfanout582 _03761_ vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__buf_2
X_16760_ clknet_leaf_28_wb_clk_i _02390_ _00456_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13972_ _03842_ _03843_ vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__nor2_1
Xfanout593 _04368_ vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__clkbuf_8
X_15711_ net1153 vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__inv_2
X_12923_ net311 net2647 net472 vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16691_ clknet_leaf_164_wb_clk_i _02321_ _00387_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08360__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13083__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15642_ net1248 vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__inv_2
X_12854_ net318 net2532 net481 vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__mux2_1
XANTENNA__11247__B1 _07104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18361_ net1346 vssd1 vssd1 vccd1 vccd1 la_data_out[9] sky130_fd_sc_hd__buf_2
X_11805_ _07616_ _07594_ _07595_ vssd1 vssd1 vccd1 vccd1 _07617_ sky130_fd_sc_hd__mux2_2
X_15573_ net1246 vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12785_ net303 net2395 net490 vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__mux2_1
X_17312_ clknet_leaf_129_wb_clk_i _02942_ _01008_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_14524_ net1063 vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__inv_2
X_11736_ _07547_ vssd1 vssd1 vccd1 vccd1 _07548_ sky130_fd_sc_hd__inv_2
X_18292_ net1384 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
XFILLER_0_84_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17243_ clknet_leaf_193_wb_clk_i _02873_ _00939_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10470__A1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14455_ net1096 vssd1 vssd1 vccd1 vccd1 _00085_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12427__S _03667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11667_ net24 net992 net918 net1937 vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__a22o_1
X_13406_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[20\]
+ net252 net416 vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__mux2_1
X_10618_ net890 _06623_ net555 vssd1 vssd1 vccd1 vccd1 _06624_ sky130_fd_sc_hd__a21o_1
X_17174_ clknet_leaf_139_wb_clk_i _02804_ _00870_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14386_ net1510 vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__clkbuf_1
X_11598_ net126 net1011 net346 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[26\]
+ vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16125_ net1136 vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__inv_2
XANTENNA__08966__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13337_ net233 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[23\]
+ net427 vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10549_ net518 _06134_ _06136_ vssd1 vssd1 vccd1 vccd1 _06559_ sky130_fd_sc_hd__and3_1
XFILLER_0_109_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16056_ net1263 vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13268_ net242 net2270 net434 vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__mux2_1
XANTENNA__12670__B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15007_ net1180 vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__inv_2
XANTENNA__13258__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08718__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12219_ _08003_ _03513_ _08004_ vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__o21a_1
XFILLER_0_110_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13199_ net243 net2302 net353 vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__mux2_1
XANTENNA__09682__D net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16958_ clknet_leaf_184_wb_clk_i _02588_ _00654_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09143__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15909_ net1288 vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16889_ clknet_leaf_12_wb_clk_i _02519_ _00585_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08351__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11506__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09430_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[5\]
+ net685 net596 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11238__B1 _07108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09361_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[7\]
+ net823 net803 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[7\]
+ _05406_ vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_19_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_74_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08312_ net944 net937 net926 vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09292_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[8\]
+ net646 net639 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[8\]
+ _05340_ vssd1 vssd1 vccd1 vccd1 _05341_ sky130_fd_sc_hd__a221o_1
XFILLER_0_118_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08243_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[31\]
+ net680 net670 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_43_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08174_ _04256_ vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10365__B _06384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08957__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput130 net130 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__buf_2
Xoutput141 net141 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__clkbuf_4
Xoutput152 net152 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__clkbuf_4
XANTENNA__13168__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08709__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout598_A net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput163 net163 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput174 net174 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__clkbuf_4
Xoutput185 net185 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__clkbuf_4
XANTENNA__12910__A0 _06499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09382__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout765_A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout386_X net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08590__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12800__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout553_X net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout932_A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14300__B team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[30\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13218__A1 _06637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09628_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[2\]
+ net700 net637 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_67_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12101__A _07864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11229__B1 _07101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_52_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09559_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[3\]
+ net715 _05592_ _05595_ vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__o22a_4
XANTENNA_fanout720_X net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout818_X net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13631__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11940__A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12570_ _03666_ net1764 net206 vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09842__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10988__C1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11521_ _07346_ _07430_ _07429_ vssd1 vssd1 vccd1 vccd1 _07432_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_156_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14240_ _04022_ _04030_ vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__nor2_1
X_11452_ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[4\] _07362_ net1002
+ vssd1 vssd1 vccd1 vccd1 _07363_ sky130_fd_sc_hd__mux2_4
XANTENNA__08026__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[24\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10403_ net896 _06420_ _05353_ vssd1 vssd1 vccd1 vccd1 _06421_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14171_ net1751 net502 net908 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[20\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__08948__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[16\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11383_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[2\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[1\]
+ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[0\] vssd1 vssd1 vccd1
+ vccd1 _07314_ sky130_fd_sc_hd__and3_1
XFILLER_0_61_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input61_A wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10334_ _05577_ _06003_ vssd1 vssd1 vccd1 vccd1 _06355_ sky130_fd_sc_hd__or2_4
X_13122_ net328 net2803 net450 vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__mux2_1
XANTENNA__08313__X _04395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13078__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17930_ clknet_leaf_43_wb_clk_i _03269_ _01626_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13053_ net304 net2463 net458 vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__mux2_1
X_10265_ _06276_ _06286_ _06288_ net537 vssd1 vssd1 vccd1 vccd1 _06289_ sky130_fd_sc_hd__a31oi_1
Xfanout1300 net1311 vssd1 vssd1 vccd1 vccd1 net1300 sky130_fd_sc_hd__buf_4
X_12004_ _07771_ _07773_ _07815_ _07658_ _07518_ vssd1 vssd1 vccd1 vccd1 _07816_ sky130_fd_sc_hd__o32a_4
Xfanout1311 net1312 vssd1 vssd1 vccd1 vccd1 net1311 sky130_fd_sc_hd__clkbuf_4
X_17861_ clknet_leaf_103_wb_clk_i _03204_ _01557_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09373__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10196_ net517 net366 _05801_ vssd1 vssd1 vccd1 vccd1 _06222_ sky130_fd_sc_hd__and3_1
XANTENNA__11180__A2 _07097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08581__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16812_ clknet_leaf_4_wb_clk_i _02442_ _00508_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17792_ clknet_leaf_92_wb_clk_i _03135_ _01488_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12710__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13457__A1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_91_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout390 _03733_ vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__buf_6
XANTENNA__09125__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16743_ clknet_leaf_203_wb_clk_i _02373_ _00439_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13955_ _03826_ _03827_ vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkload7_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12906_ net254 net2188 net472 vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__mux2_1
XANTENNA__11553__C _07434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16674_ clknet_leaf_8_wb_clk_i _02304_ _00370_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13886_ net1596 net982 _03779_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[14\]
+ sky130_fd_sc_hd__o21a_1
X_18413_ net183 vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15625_ net1159 vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12837_ net230 net2147 net481 vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13541__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18344_ net1333 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
XFILLER_0_16_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15556_ net1117 vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__inv_2
X_12768_ net234 net2402 net490 vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__mux2_1
XANTENNA__09833__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18355__1340 vssd1 vssd1 vccd1 vccd1 _18355__1340/HI net1340 sky130_fd_sc_hd__conb_1
XANTENNA__12665__B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10737__Y _06737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14507_ net1067 vssd1 vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__inv_2
X_18275_ clknet_leaf_37_wb_clk_i _03504_ _01970_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[29\]
+ sky130_fd_sc_hd__dfrtp_4
X_11719_ _07519_ _07530_ vssd1 vssd1 vccd1 vccd1 _07531_ sky130_fd_sc_hd__nand2_1
X_15487_ net1156 vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__inv_2
X_12699_ net238 net2391 net498 vssd1 vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__mux2_1
XANTENNA__10994__A2 _06540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09677__D net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17226_ clknet_leaf_196_wb_clk_i _02856_ _00922_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_14438_ net1280 vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__inv_2
Xinput10 DAT_I[17] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput21 DAT_I[27] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
Xinput32 DAT_I[8] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
Xinput43 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__clkbuf_1
Xinput54 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08939__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17157_ clknet_leaf_176_wb_clk_i _02787_ _00853_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput65 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_1
Xhold805 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[12\] vssd1
+ vssd1 vccd1 vccd1 net2219 sky130_fd_sc_hd__dlygate4sd3_1
X_14369_ _04128_ _04141_ _04123_ vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__o21ai_1
Xhold816 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2230 sky130_fd_sc_hd__dlygate4sd3_1
X_16108_ net1308 vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold827 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2241 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_137_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_137_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold838 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net2252 sky130_fd_sc_hd__dlygate4sd3_1
Xhold849 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2263 sky130_fd_sc_hd__dlygate4sd3_1
X_17088_ clknet_leaf_130_wb_clk_i _02718_ _00784_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08930_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[16\]
+ net822 net737 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04994_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16039_ net1284 vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09990__A _05256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09364__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08861_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[17\]
+ net663 net611 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__a22o_1
XANTENNA__17980__Q net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11171__A2 _07117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08572__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1505 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net2919 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1516 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2930 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12620__S _03682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08792_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[19\]
+ net814 net806 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__a22o_1
Xhold1527 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 net2941 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1538 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 net2952 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1549 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2963 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09116__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_918 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09413_ _05451_ _05453_ _05455_ _05456_ vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__or4_1
XANTENNA__13451__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1088_A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09344_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[7\]
+ net666 net661 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[7\]
+ _05390_ vssd1 vssd1 vccd1 vccd1 _05391_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09824__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09275_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[9\]
+ net827 net784 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_136_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout513_A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1255_A net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08226_ net884 net869 net858 vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09037__D1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08157_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[4\] team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_151_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1092 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08088_ net1025 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[17\]
+ net971 _04193_ vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18400__1372 vssd1 vssd1 vccd1 vccd1 _18400__1372/HI net1372 sky130_fd_sc_hd__conb_1
XANTENNA__09355__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10050_ _06077_ _06078_ vssd1 vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout670_X net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08787__Y _04858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08563__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout768_X net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13626__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12530__S net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12102__Y _07914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout935_X net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08315__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13740_ net923 _06623_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[8\]
+ sky130_fd_sc_hd__nor2_1
X_10952_ net961 _06387_ net567 vssd1 vssd1 vccd1 vccd1 _06939_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_175_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13671_ net2619 net257 net384 vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__mux2_1
X_10883_ _06787_ _06879_ _06784_ _06785_ vssd1 vssd1 vccd1 vccd1 _06880_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_123_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11670__A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15410_ net1140 vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__inv_2
XFILLER_0_168_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12622_ _03655_ net1803 net202 vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__mux2_1
X_16390_ clknet_leaf_119_wb_clk_i _02020_ _00086_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09815__B1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13611__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15341_ net1082 vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12553_ _03646_ net2096 net207 vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__mux2_1
XANTENNA__08094__A2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[14\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18060_ net1037 _03398_ _01756_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[15\]
+ sky130_fd_sc_hd__dfrtp_4
X_11504_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[10\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[10\]
+ net1034 vssd1 vssd1 vccd1 vccd1 _07415_ sky130_fd_sc_hd__mux2_1
X_15272_ net1223 vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__inv_2
X_12484_ net1696 _03646_ net210 vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17011_ clknet_leaf_164_wb_clk_i _02641_ _00707_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_14223_ team_05_WB.instance_to_wrap.total_design.keypad0.counter\[3\] team_05_WB.instance_to_wrap.total_design.keypad0.counter\[4\]
+ team_05_WB.instance_to_wrap.total_design.keypad0.counter\[5\] _04017_ vssd1 vssd1
+ vccd1 vccd1 _04019_ sky130_fd_sc_hd__and4_1
X_11435_ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[31\] _07347_ net1003
+ vssd1 vssd1 vccd1 vccd1 _07348_ sky130_fd_sc_hd__mux2_1
XANTENNA__13914__A2 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10189__B1 _06215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12705__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1012 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11366_ _07305_ team_05_WB.instance_to_wrap.total_design.data_from_keypad\[0\] net509
+ vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__mux2_1
X_14154_ _03838_ net907 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[3\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__09594__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10317_ net338 _06333_ _06338_ net336 vssd1 vssd1 vccd1 vccd1 _06339_ sky130_fd_sc_hd__o22a_1
X_13105_ net246 net2798 net450 vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11548__C _07394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11297_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[73\] _07109_
+ _07113_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[41\] _07214_
+ vssd1 vssd1 vccd1 vccd1 _07257_ sky130_fd_sc_hd__a221o_1
X_14085_ _03950_ _03951_ vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08203__B net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09346__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17913_ clknet_leaf_99_wb_clk_i _03256_ _01609_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10248_ _04637_ _04678_ _05906_ vssd1 vssd1 vccd1 vccd1 _06272_ sky130_fd_sc_hd__or3_1
X_13036_ net237 net2518 net459 vssd1 vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__mux2_1
Xfanout1130 net1137 vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__clkbuf_2
Xfanout1141 net1151 vssd1 vssd1 vccd1 vccd1 net1141 sky130_fd_sc_hd__buf_2
XANTENNA__11845__A team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13536__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17844_ clknet_leaf_88_wb_clk_i _03187_ _01540_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[90\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1152 net1153 vssd1 vssd1 vccd1 vccd1 net1152 sky130_fd_sc_hd__buf_4
X_10179_ _06008_ _06015_ net516 vssd1 vssd1 vccd1 vccd1 _06206_ sky130_fd_sc_hd__mux2_1
Xfanout1163 net1177 vssd1 vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__clkbuf_4
Xfanout1174 net1175 vssd1 vssd1 vccd1 vccd1 net1174 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10900__A2 _06108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1185 net1186 vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__buf_2
XFILLER_0_89_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17775_ clknet_leaf_89_wb_clk_i _03118_ _01471_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1196 net1198 vssd1 vssd1 vccd1 vccd1 net1196 sky130_fd_sc_hd__buf_4
X_14987_ net1077 vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10113__A0 _06125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16726_ clknet_leaf_140_wb_clk_i _02356_ _00422_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13938_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[5\] team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__or2_1
XFILLER_0_135_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16657_ clknet_leaf_169_wb_clk_i _02287_ _00353_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13869_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[6\]
+ net559 net575 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[6\]
+ net986 vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13271__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15608_ net1168 vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16588_ clknet_leaf_0_wb_clk_i _02218_ _00284_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08218__X _04301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10467__Y _06481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18327_ net1318 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
XANTENNA__10416__A1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15539_ net1140 vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_40_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09060_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[13\]
+ net679 net628 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[13\]
+ _05107_ vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__a221o_1
X_18258_ clknet_leaf_39_wb_clk_i _03487_ _01953_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09985__A net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17209_ clknet_leaf_15_wb_clk_i _02839_ _00905_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12615__S net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18189_ clknet_leaf_42_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[10\]
+ _01884_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_163_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold602 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 net2016 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold613 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 net2027 sky130_fd_sc_hd__dlygate4sd3_1
Xhold624 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2038 sky130_fd_sc_hd__dlygate4sd3_1
Xhold635 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2049 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold646 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net2060 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08793__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold657 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2071 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold668 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2082 sky130_fd_sc_hd__dlygate4sd3_1
X_09962_ _05902_ _05990_ vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__nand2_1
Xhold679 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net2093 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08913_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[16\]
+ net672 net644 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__a22o_1
XANTENNA__09337__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09893_ net891 _05921_ vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13446__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08545__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1302 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net2716 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08844_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[18\]
+ net837 net752 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[18\]
+ _04911_ vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__a221o_1
Xhold1313 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net2727 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1003_A _07345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10649__A2_N net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1324 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1335 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2749 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1346 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 net2760 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1357 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2771 sky130_fd_sc_hd__dlygate4sd3_1
X_08775_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[19\]
+ net680 net630 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[19\]
+ _04845_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__a221o_1
Xhold1368 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2782 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout463_A _03711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold1379 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net2793 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10655__A1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout630_A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout728_A net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11490__A _07346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13181__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09327_ net572 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[8\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[8\] vssd1 vssd1 vccd1
+ vccd1 _05374_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11604__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09258_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[29\] _05308_
+ vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_170_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08209_ net884 net869 net864 vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__and3_4
XFILLER_0_90_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12525__S net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09189_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[10\]
+ net711 net672 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[10\]
+ _05241_ vssd1 vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11220_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[61\] _07115_
+ _07117_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[53\] _07183_
+ vssd1 vssd1 vccd1 vccd1 _07184_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_79_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13109__A0 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout885_X net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08784__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11151_ _07060_ _07112_ vssd1 vssd1 vccd1 vccd1 _07117_ sky130_fd_sc_hd__nor2_4
XANTENNA__10591__B1 _06284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10102_ net375 net361 vssd1 vssd1 vccd1 vccd1 _06130_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11082_ _04162_ _04163_ _07041_ vssd1 vssd1 vccd1 vccd1 _07049_ sky130_fd_sc_hd__or3b_1
XANTENNA__13356__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10033_ _05531_ _06061_ vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__nor2_1
X_14910_ net1054 vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__inv_2
X_15890_ net1296 vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__inv_2
XANTENNA_input24_A DAT_I[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14841_ net1053 vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_125_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17560_ clknet_leaf_59_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[31\]
+ _01256_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_14772_ net1066 vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__inv_2
X_11984_ _07777_ _07786_ _07795_ net356 vssd1 vssd1 vccd1 vccd1 _07796_ sky130_fd_sc_hd__o31a_4
XFILLER_0_169_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16511_ clknet_leaf_156_wb_clk_i _02141_ _00207_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13723_ net905 _06350_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[23\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__09500__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10935_ net1043 _06923_ _06924_ net960 vssd1 vssd1 vccd1 vccd1 _06925_ sky130_fd_sc_hd__a211o_1
X_17491_ clknet_leaf_36_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[26\]
+ _01187_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13091__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16442_ clknet_leaf_31_wb_clk_i _02072_ _00138_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13654_ net2571 net310 net388 vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10866_ _06812_ _06862_ vssd1 vssd1 vccd1 vccd1 _06863_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12399__A1 _07816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12605_ net1635 _07821_ _03680_ vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16373_ clknet_leaf_175_wb_clk_i _02003_ _00069_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13585_ net2125 net317 net396 vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__mux2_1
X_10797_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[22\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06794_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18112_ clknet_leaf_69_wb_clk_i _03435_ _01808_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[29\]
+ sky130_fd_sc_hd__dfstp_2
X_15324_ net1064 vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__inv_2
X_12536_ _07821_ net1909 _03675_ vssd1 vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18043_ clknet_leaf_54_wb_clk_i _03381_ _01739_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_30_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15255_ net1097 vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__inv_2
X_12467_ net1730 _07821_ _03670_ vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__mux2_1
XANTENNA__12435__S _03667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14206_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[9\] _04006_
+ vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_144_Right_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11418_ _07324_ _07338_ vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15186_ net1233 vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__inv_2
X_12398_ net1769 _07821_ _07852_ vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__mux2_1
XANTENNA__08214__A net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12571__A1 _07821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08775__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14137_ net1751 net502 net911 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[20\]
+ sky130_fd_sc_hd__and3_1
X_11349_ net980 net508 _07296_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14068_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[11\] _03884_ vssd1
+ vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__nand2_1
XANTENNA__08527__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13266__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13019_ net294 net2271 net463 vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17827_ clknet_leaf_87_wb_clk_i _03170_ _01523_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[73\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08560_ _04634_ _04635_ vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__or2_1
X_17758_ clknet_leaf_84_wb_clk_i _03101_ _01454_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10637__A1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08491_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[27\]
+ net653 net618 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__a22o_1
X_16709_ clknet_leaf_179_wb_clk_i _02339_ _00405_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17689_ clknet_leaf_99_wb_clk_i _03032_ _01385_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[127\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11514__S net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09112_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[12\]
+ net767 net748 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_152_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_152_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09043_ _05078_ _05100_ vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__and2_2
XFILLER_0_4_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout211_A _03674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold410 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[26\] vssd1 vssd1
+ vccd1 vccd1 net1824 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold421 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[49\] vssd1 vssd1
+ vccd1 vccd1 net1835 sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[103\] vssd1 vssd1
+ vccd1 vccd1 net1846 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12562__A1 _07812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold443 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[95\] vssd1 vssd1
+ vccd1 vccd1 net1857 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold454 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[50\] vssd1 vssd1
+ vccd1 vccd1 net1868 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1120_A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold465 net135 vssd1 vssd1 vccd1 vccd1 net1879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 team_05_WB.instance_to_wrap.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 net1890
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold487 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[33\] vssd1 vssd1
+ vccd1 vccd1 net1901 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout901 net902 vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__clkbuf_2
Xhold498 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1912 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout912 _03797_ vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__buf_2
X_09945_ _05932_ _05973_ _05931_ vssd1 vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__a21oi_1
Xfanout923 _05213_ vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout580_A net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout934 _04372_ vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13176__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08518__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout678_A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout945 _04364_ vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__buf_2
Xfanout956 net958 vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ _05904_ vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__inv_2
Xfanout967 net968 vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__buf_2
Xhold1110 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[8\] vssd1 vssd1
+ vccd1 vccd1 net2524 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout978 team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[14\] vssd1 vssd1
+ vccd1 vccd1 net978 sky130_fd_sc_hd__buf_2
Xfanout989 _07482_ vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__buf_2
Xhold1121 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2535 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09191__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1132 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2546 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ _04889_ _04891_ _04893_ _04895_ vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__or4_1
XANTENNA__09730__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1143 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 net2557 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout845_A _04373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout466_X net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1154 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 net2568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1165 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net2579 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1176 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2590 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1187 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net2601 sky130_fd_sc_hd__dlygate4sd3_1
X_08758_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[21\]
+ net851 _04827_ _04829_ net855 vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__a2111o_1
Xhold1198 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 net2612 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08297__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08689_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[22\]
+ net704 net658 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout633_X net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10720_ net2377 net309 net539 vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_172_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10651_ net1991 net303 net540 vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout800_X net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11053__A1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10582_ _05958_ _06589_ vssd1 vssd1 vccd1 vccd1 _06590_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13370_ net2158 net230 net422 vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12321_ net547 net354 vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__nand2_4
XFILLER_0_133_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09549__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15040_ net1198 vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__inv_2
X_12252_ _03545_ _03546_ _03511_ vssd1 vssd1 vccd1 vccd1 _03547_ sky130_fd_sc_hd__o21a_1
XFILLER_0_107_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08757__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11203_ net149 net731 _07160_ _07167_ vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__o22a_1
XANTENNA__17345__CLK clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12183_ _07991_ _07992_ _07988_ _07989_ vssd1 vssd1 vccd1 vccd1 _07995_ sky130_fd_sc_hd__a2bb2o_1
X_11134_ _07087_ _07098_ vssd1 vssd1 vccd1 vccd1 _07100_ sky130_fd_sc_hd__nor2_4
X_16991_ clknet_leaf_153_wb_clk_i _02621_ _00687_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13086__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11065_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[2\] team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[1\]
+ vssd1 vssd1 vccd1 vccd1 _07032_ sky130_fd_sc_hd__or2_1
X_15942_ net1272 vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__inv_2
XANTENNA__09182__B1 _05215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10016_ _06043_ _06044_ vssd1 vssd1 vccd1 vccd1 _06045_ sky130_fd_sc_hd__nand2_1
X_15873_ net1269 vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__inv_2
X_17612_ clknet_leaf_57_wb_clk_i _02983_ _01308_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_14824_ net1219 vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__inv_2
X_17543_ clknet_leaf_61_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[14\]
+ _01239_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10619__A1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14755_ net1203 vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11967_ _07726_ _07743_ vssd1 vssd1 vccd1 vccd1 _07779_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_59_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13706_ net900 _06658_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[6\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_80_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10918_ net961 _06910_ vssd1 vssd1 vccd1 vccd1 _06911_ sky130_fd_sc_hd__or2_1
X_17474_ clknet_leaf_41_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[9\]
+ _01170_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14686_ net1054 vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11898_ _07685_ _07686_ _07707_ _07708_ vssd1 vssd1 vccd1 vccd1 _07710_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16425_ clknet_leaf_18_wb_clk_i _02055_ _00121_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13637_ net2222 net254 net388 vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10849_ _06835_ _06836_ _06845_ vssd1 vssd1 vccd1 vccd1 _06846_ sky130_fd_sc_hd__and3_1
XFILLER_0_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11044__A1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10666__A1_N team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16356_ clknet_leaf_179_wb_clk_i _01986_ _00052_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13568_ net2300 net232 net398 vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__mux2_1
XANTENNA__12673__B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10252__C1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15307_ net1071 vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12519_ net1743 _03655_ net208 vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__mux2_1
X_16287_ net1253 vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13499_ net2483 net244 net406 vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__mux2_1
XANTENNA__08460__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09685__D net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18026_ clknet_leaf_97_wb_clk_i _03365_ _01722_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_wire381_A _04342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15238_ net1208 vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08748__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_2_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15169_ net1224 vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout208 _03676_ vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__buf_4
XANTENNA__08231__X _04314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout219 net221 vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10480__Y _06494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_52_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09730_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[0\]
+ net795 _05741_ _05747_ _05754_ vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_157_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09661_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[1\]
+ net781 _05674_ _05675_ _05686_ vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__a2111oi_1
XTAP_TAPCELL_ROW_2_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08920__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08612_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[24\]
+ net693 net661 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__a22o_1
X_09592_ _05624_ _05625_ _05626_ _05627_ vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_141_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08543_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[26\]
+ net758 net747 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[26\]
+ _04618_ vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__a221o_1
XFILLER_0_82_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout259_A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10086__A2 _05801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08474_ _04552_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[28\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_9_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout426_A _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1168_A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08987__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout214_X net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08451__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09026_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[14\]
+ net839 net757 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[14\]
+ _05085_ vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_76_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12535__A1 _03666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08739__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout795_A _04395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold240 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[11\] vssd1 vssd1
+ vccd1 vccd1 net1654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[80\] vssd1 vssd1
+ vccd1 vccd1 net1665 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12803__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09400__B2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[26\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold262 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[26\]
+ vssd1 vssd1 vccd1 vccd1 net1676 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 team_05_WB.instance_to_wrap.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 net1687
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold284 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[94\] vssd1 vssd1
+ vccd1 vccd1 net1698 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[99\] vssd1 vssd1
+ vccd1 vccd1 net1709 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10390__Y _06408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout962_A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout720 _04285_ vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14303__B _04552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout731 _07030_ vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_165_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09928_ net349 _05330_ _05378_ _05955_ _05939_ vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__o221ai_4
Xfanout742 net744 vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__clkbuf_8
Xfanout753 net755 vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__buf_6
Xfanout764 net767 vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09164__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08301__B net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout775 net777 vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__buf_6
Xfanout786 _04400_ vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__clkbuf_8
X_09859_ _04879_ _05840_ _05884_ _05887_ _04881_ vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__a2111o_2
XANTENNA_fanout750_X net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout797 _04395_ vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_172_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout848_X net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08911__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13634__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12870_ net230 net2113 net478 vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__mux2_1
X_11821_ _07621_ _07625_ _07627_ _07630_ _07631_ vssd1 vssd1 vccd1 vccd1 _07633_ sky130_fd_sc_hd__a2111o_2
XANTENNA__10559__A net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10077__A2 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14540_ net1072 vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__inv_2
X_11752_ _07554_ _07557_ vssd1 vssd1 vccd1 vccd1 _07564_ sky130_fd_sc_hd__nand2b_1
XANTENNA__08029__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[20\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10703_ _06701_ _06704_ _04264_ vssd1 vssd1 vccd1 vccd1 _06705_ sky130_fd_sc_hd__a21oi_4
X_14471_ net1105 vssd1 vssd1 vccd1 vccd1 _00101_ sky130_fd_sc_hd__inv_2
X_11683_ net43 net42 net45 net44 vssd1 vssd1 vccd1 vccd1 _07497_ sky130_fd_sc_hd__or4_1
XANTENNA__14318__X _04091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08690__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16210_ net1212 vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__inv_2
XANTENNA__11026__A1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13422_ net2286 net328 net418 vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__mux2_1
X_10634_ _05423_ _05954_ vssd1 vssd1 vccd1 vccd1 _06639_ sky130_fd_sc_hd__xor2_1
XANTENNA__08427__C1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17190_ clknet_leaf_116_wb_clk_i _02820_ _00886_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16141_ net1274 vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08978__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13353_ net304 net2851 net426 vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10565_ _05826_ _05959_ vssd1 vssd1 vccd1 vccd1 _06574_ sky130_fd_sc_hd__nand2_1
XANTENNA__08442__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12304_ _03511_ _03557_ _03569_ _03575_ vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__and4_1
X_16072_ net1169 vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13284_ net286 net2308 net432 vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__mux2_1
X_10496_ net369 net347 vssd1 vssd1 vccd1 vccd1 _06509_ sky130_fd_sc_hd__nor2_1
XANTENNA__12526__A1 _03645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15023_ net1233 vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__inv_2
X_12235_ _03511_ _03524_ _03528_ _03529_ _07992_ vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__a32oi_4
XANTENNA__12713__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12166_ _07968_ _07977_ vssd1 vssd1 vccd1 vccd1 _07978_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_9_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11117_ _07072_ _07083_ vssd1 vssd1 vccd1 vccd1 _07084_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16974_ clknet_leaf_171_wb_clk_i _02604_ _00670_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_12097_ _07908_ vssd1 vssd1 vccd1 vccd1 _07909_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_30_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15925_ net1256 vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__inv_2
X_11048_ _04170_ _06085_ _06718_ _07016_ net960 vssd1 vssd1 vccd1 vccd1 _07017_ sky130_fd_sc_hd__a311o_1
Xinput8 DAT_I[15] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XANTENNA__13544__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15856_ net1273 vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__inv_2
XANTENNA__12668__B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14807_ net1099 vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__inv_2
X_15787_ net1301 vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__inv_2
XANTENNA__10469__A net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12999_ net218 net2505 net463 vssd1 vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14738_ net1238 vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__inv_2
X_17526_ clknet_leaf_113_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[29\]
+ _01222_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_157_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17457_ clknet_leaf_65_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[25\]
+ _01153_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14375__S _00040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14669_ net1080 vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08681__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16408_ clknet_leaf_30_wb_clk_i _02038_ _00104_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_08190_ net1019 _04272_ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__nand2_1
X_17388_ clknet_leaf_58_wb_clk_i net1448 _01084_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11568__A2 _07354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08969__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16339_ net1125 vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09993__A _05350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_144_Left_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18009_ clknet_leaf_63_wb_clk_i _03348_ _01705_ vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12623__S net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09394__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10370__C _05978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09146__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09713_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[0\]
+ net1017 net944 net926 vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__and4_1
XANTENNA__13454__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09644_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[1\]
+ net946 net1013 net924 vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_153_Left_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09575_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[2\]
+ net941 net1013 net924 vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__and4_1
XFILLER_0_139_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_42_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08526_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[26\]
+ net616 net612 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__a22o_1
XANTENNA__08657__C1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08457_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[28\]
+ net817 net807 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__a22o_1
XANTENNA__08672__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout429_X net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout808_A net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08388_ _04467_ vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08424__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18281__A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_162_Left_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10350_ net893 _06369_ vssd1 vssd1 vccd1 vccd1 _06370_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_115_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout798_X net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13629__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09009_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[14\]
+ net708 net678 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10281_ net531 _06191_ net333 vssd1 vssd1 vccd1 vccd1 _06304_ sky130_fd_sc_hd__a21o_1
XANTENNA__12533__S net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13856__C net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14314__A net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12020_ _07816_ _07819_ _07821_ _07831_ vssd1 vssd1 vccd1 vccd1 _07832_ sky130_fd_sc_hd__and4_1
XANTENNA__09385__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11192__B1 _07101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10561__B _06570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08312__A net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout550 _07448_ vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09137__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_81_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout561 team_05_WB.instance_to_wrap.total_design.core.data_mem.next_write vssd1
+ vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__buf_2
Xfanout572 net573 vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__buf_2
X_13971_ _03821_ _03840_ _03841_ vssd1 vssd1 vccd1 vccd1 _03843_ sky130_fd_sc_hd__nor3_1
Xfanout594 net597 vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__buf_6
XPHY_EDGE_ROW_171_Left_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15710_ net1165 vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__inv_2
XANTENNA__13364__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12922_ net330 net2434 net474 vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__mux2_1
X_16690_ clknet_leaf_127_wb_clk_i _02320_ _00386_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15641_ net1250 vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__inv_2
X_12853_ net303 net2170 net482 vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18360_ net1345 vssd1 vssd1 vccd1 vccd1 la_data_out[8] sky130_fd_sc_hd__buf_2
X_11804_ _07580_ _07594_ vssd1 vssd1 vccd1 vccd1 _07616_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15572_ net1282 vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__inv_2
X_12784_ net295 net2860 net491 vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17311_ clknet_leaf_152_wb_clk_i _02941_ _01007_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_84_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14523_ net1098 vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__inv_2
X_11735_ _07540_ _07546_ _07533_ vssd1 vssd1 vccd1 vccd1 _07547_ sky130_fd_sc_hd__o21a_2
X_18291_ net1383 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
XANTENNA__12708__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08663__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17242_ clknet_leaf_10_wb_clk_i _02872_ _00938_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14454_ net1084 vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__inv_2
XANTENNA__10470__A2 _06481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11666_ net27 net992 _07483_ net2104 vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13405_ net2504 net246 net418 vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__mux2_1
X_10617_ _05378_ _05815_ vssd1 vssd1 vccd1 vccd1 _06623_ sky130_fd_sc_hd__xnor2_2
X_17173_ clknet_leaf_175_wb_clk_i _02803_ _00869_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_14385_ net1518 vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08415__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11597_ net1682 net1009 net345 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[27\]
+ vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16124_ net1136 vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__inv_2
X_13336_ net235 net2607 net427 vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__mux2_1
X_10548_ _06556_ _06557_ net889 vssd1 vssd1 vccd1 vccd1 _06558_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13539__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16055_ net1262 vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__inv_2
XANTENNA__12443__S net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13267_ net222 net2364 net434 vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10479_ net554 _06484_ _06492_ net348 vssd1 vssd1 vccd1 vccd1 _06493_ sky130_fd_sc_hd__o22a_1
X_15006_ net1056 vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__inv_2
X_12218_ _08000_ _08006_ vssd1 vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__nor2_1
XANTENNA__09950__A_N _04818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13198_ _06270_ net2668 net352 vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__mux2_1
XANTENNA__10471__B net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12149_ _07911_ _07950_ _07958_ vssd1 vssd1 vccd1 vccd1 _07961_ sky130_fd_sc_hd__and3b_1
XANTENNA__10930__B1 _06898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16957_ clknet_leaf_128_wb_clk_i _02587_ _00653_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13274__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15908_ net1296 vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16888_ clknet_leaf_33_wb_clk_i _02518_ _00584_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15839_ net1292 vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09360_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[7\]
+ net847 net734 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_802 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08311_ net948 net937 net925 vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__and3_1
X_17509_ clknet_leaf_74_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[12\]
+ _01205_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_09291_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[8\]
+ net705 net702 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__a22o_1
XANTENNA__12618__S _03682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08654__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11522__S net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_126_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_118_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1081 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08242_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[31\]
+ net653 net638 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_59_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_16_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08173_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[10\] team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[9\]
+ _04249_ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__and3_1
XANTENNA__08406__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13449__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput120 net120 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__buf_2
Xoutput131 net131 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1033_A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xoutput142 net142 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__clkbuf_4
XANTENNA__09367__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput153 net153 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__clkbuf_4
XANTENNA__09228__A net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput164 net164 vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_110_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput175 net175 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__clkbuf_4
XANTENNA__11174__B1 _07130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout493_A _03699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput186 net186 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__clkbuf_4
XANTENNA__09119__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout660_A net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13184__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout758_A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11493__A _07346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_165_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09627_ _05658_ _05659_ _05660_ _05661_ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_108_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13218__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout546_X net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08893__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout925_A net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12426__A0 _03604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09558_ _05582_ _05583_ _05585_ _05594_ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__or4_1
XFILLER_0_84_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08509_ _04580_ _04582_ _04584_ _04586_ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__or4_1
XFILLER_0_77_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12528__S _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09489_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[4\]
+ net851 net847 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[4\]
+ _05518_ vssd1 vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__a221o_1
XANTENNA__08645__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout713_X net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11520_ _07346_ _07430_ _07429_ vssd1 vssd1 vccd1 vccd1 _07431_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_156_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11451_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[4\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[4\]
+ net1035 vssd1 vssd1 vccd1 vccd1 _07362_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10402_ _06097_ _06419_ vssd1 vssd1 vccd1 vccd1 _06420_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14170_ net2306 net503 net909 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[19\]
+ sky130_fd_sc_hd__and3_1
X_11382_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[1\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[0\]
+ vssd1 vssd1 vccd1 vccd1 _07313_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09070__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13359__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13121_ net314 net2781 net451 vssd1 vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__mux2_1
X_10333_ net1021 _04756_ _04757_ net552 vssd1 vssd1 vccd1 vccd1 _06354_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09358__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input54_A wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13052_ net295 net2913 net458 vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__mux2_1
X_10264_ _05577_ _06049_ _06287_ net510 _04636_ vssd1 vssd1 vccd1 vccd1 _06288_ sky130_fd_sc_hd__o32a_1
XANTENNA__11165__B1 _07109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12003_ _07765_ _07767_ _07769_ vssd1 vssd1 vccd1 vccd1 _07815_ sky130_fd_sc_hd__nor3_1
Xfanout1301 net1303 vssd1 vssd1 vccd1 vccd1 net1301 sky130_fd_sc_hd__buf_4
Xfanout1312 net1313 vssd1 vssd1 vccd1 vccd1 net1312 sky130_fd_sc_hd__buf_4
X_17860_ clknet_leaf_80_wb_clk_i _03203_ _01556_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[42\]
+ sky130_fd_sc_hd__dfrtp_1
X_10195_ net893 _06218_ _06220_ net556 vssd1 vssd1 vccd1 vccd1 _06221_ sky130_fd_sc_hd__a211o_1
X_16811_ clknet_leaf_188_wb_clk_i _02441_ _00507_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_17791_ clknet_leaf_89_wb_clk_i _03134_ _01487_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[101\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout391 _03733_ vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__buf_4
X_13954_ net980 _03812_ _03813_ vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__a21boi_1
X_16742_ clknet_leaf_116_wb_clk_i _02372_ _00438_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09530__B1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12905_ net249 net2722 net474 vssd1 vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__mux2_1
X_16673_ clknet_leaf_147_wb_clk_i _02303_ _00369_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13885_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[14\]
+ net560 net576 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[14\]
+ net987 vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__a221o_1
XANTENNA__08884__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11690__X net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12417__A0 _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18412_ net1376 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__buf_2
XFILLER_0_69_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15624_ net1160 vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12836_ net234 net2899 net481 vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__mux2_1
XANTENNA__09160__X _05215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18343_ net1332 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
X_15555_ net1131 vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1087 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12767_ net240 net2561 net490 vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08636__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14506_ net1116 vssd1 vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__inv_2
XFILLER_0_166_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18274_ clknet_leaf_38_wb_clk_i _03503_ _01969_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[28\]
+ sky130_fd_sc_hd__dfrtp_4
X_11718_ _07379_ _07447_ _07524_ vssd1 vssd1 vccd1 vccd1 _07530_ sky130_fd_sc_hd__or3_2
XFILLER_0_166_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15486_ net1154 vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12698_ net243 net2761 net498 vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14437_ net1191 vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17225_ clknet_leaf_21_wb_clk_i _02855_ _00921_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput11 DAT_I[18] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
X_11649_ net14 net989 net916 net1751 vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__o22a_1
XFILLER_0_86_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput22 DAT_I[28] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput33 DAT_I[9] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
Xinput44 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17156_ clknet_leaf_186_wb_clk_i _02786_ _00852_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput55 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
X_14368_ _04136_ _04140_ _04082_ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__a21oi_1
Xinput66 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09061__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12681__B net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold806 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2220 sky130_fd_sc_hd__dlygate4sd3_1
X_16107_ net1310 vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__inv_2
Xhold817 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2231 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13269__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13319_ net2005 net294 net430 vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__mux2_1
Xhold828 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2242 sky130_fd_sc_hd__dlygate4sd3_1
X_17087_ clknet_leaf_153_wb_clk_i _02717_ _00783_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold839 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 net2253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14299_ _04490_ _04510_ vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16038_ net1243 vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_177_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_177_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08860_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[17\]
+ net686 net637 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__a22o_1
XANTENNA__12901__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1506 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2920 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_106_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_106_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold1517 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2931 sky130_fd_sc_hd__dlygate4sd3_1
X_08791_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[19\]
+ net772 net746 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[19\]
+ _04860_ vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__a221o_1
X_17989_ clknet_leaf_83_wb_clk_i _03328_ _01685_ vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__dfrtp_1
Xhold1528 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2942 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1539 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2953 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12656__B1 team_05_WB.instance_to_wrap.total_design.core.instr_fetch vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09521__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08875__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12408__A0 _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09412_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[6\]
+ net850 net733 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[6\]
+ _05445_ vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__a221o_1
XANTENNA__15513__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09343_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[7\]
+ net626 net612 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__a22o_1
XANTENNA__08627__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17501__Q team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_158_Right_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout339_A _03693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09230__B _05256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09274_ _05317_ _05319_ _05321_ _05323_ vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_134_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08225_ net883 net867 net862 vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1150_A net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout506_A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1248_A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08156_ _04231_ net1022 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__or3b_2
XFILLER_0_99_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_151_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09052__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13179__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08087_ net1025 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__and2b_1
XFILLER_0_28_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1036_X net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout496_X net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12811__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input1_X net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08989_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[15\]
+ net802 net737 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[15\]
+ _05050_ vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout663_X net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_127_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10951_ _06935_ _06936_ _06937_ net961 vssd1 vssd1 vccd1 vccd1 _06938_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout830_X net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08866__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13642__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13670_ net2176 net254 net384 vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10882_ _06786_ _06878_ vssd1 vssd1 vccd1 vccd1 _06879_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_123_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11670__B team_05_WB.instance_to_wrap.total_design.core.instr_fetch vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12621_ _03646_ net1878 _03683_ vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__mux2_1
XANTENNA__09421__A _05442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08618__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15340_ net1072 vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__inv_2
X_12552_ net1738 _07793_ _03678_ vssd1 vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09291__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18317__1409 vssd1 vssd1 vccd1 vccd1 net1409 _18317__1409/LO sky130_fd_sc_hd__conb_1
XFILLER_0_53_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11503_ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[19\] _07413_ net1003
+ vssd1 vssd1 vccd1 vccd1 _07414_ sky130_fd_sc_hd__mux2_2
XFILLER_0_53_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15271_ net1106 vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__inv_2
X_12483_ net1718 _07793_ _03673_ vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__mux2_1
X_17010_ clknet_leaf_123_wb_clk_i _02640_ _00706_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_14222_ team_05_WB.instance_to_wrap.total_design.keypad0.counter\[3\] _04017_ vssd1
+ vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11434_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[31\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[31\]
+ net1033 vssd1 vssd1 vccd1 vccd1 _07347_ sky130_fd_sc_hd__mux2_1
XANTENNA__10189__A1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08324__X _04406_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12104__A_N _07914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13089__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14153_ _03820_ _03994_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[2\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11365_ _07286_ _07291_ _07293_ _07299_ _07304_ vssd1 vssd1 vccd1 vccd1 _07305_ sky130_fd_sc_hd__a311o_1
XANTENNA__08251__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10506__S net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_4_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13104_ net229 net2425 net451 vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__mux2_1
XANTENNA__14324__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10316_ _06337_ vssd1 vssd1 vccd1 vccd1 _06338_ sky130_fd_sc_hd__inv_2
X_14084_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[10\] net979 team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__a21o_1
X_11296_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[57\] _07115_
+ _07117_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[49\] _07255_
+ vssd1 vssd1 vccd1 vccd1 _07256_ sky130_fd_sc_hd__a221o_1
X_17912_ clknet_leaf_104_wb_clk_i _03255_ _01608_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13035_ net240 net2694 net458 vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__mux2_1
XANTENNA__12721__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10247_ net2201 net223 net540 vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__mux2_1
Xfanout1120 net1127 vssd1 vssd1 vccd1 vccd1 net1120 sky130_fd_sc_hd__clkbuf_2
Xfanout1131 net1133 vssd1 vssd1 vccd1 vccd1 net1131 sky130_fd_sc_hd__buf_4
XANTENNA__12350__A2 _07476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1142 net1151 vssd1 vssd1 vccd1 vccd1 net1142 sky130_fd_sc_hd__buf_4
X_17843_ clknet_leaf_90_wb_clk_i _03186_ _01539_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[89\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1153 net1163 vssd1 vssd1 vccd1 vccd1 net1153 sky130_fd_sc_hd__buf_4
X_10178_ net512 _06005_ vssd1 vssd1 vccd1 vccd1 _06205_ sky130_fd_sc_hd__or2_1
Xfanout1164 net1165 vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__buf_4
Xfanout1175 net1177 vssd1 vssd1 vccd1 vccd1 net1175 sky130_fd_sc_hd__buf_2
XANTENNA__12638__A0 _03666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1186 net1211 vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__clkbuf_2
X_17774_ clknet_leaf_87_wb_clk_i _03117_ _01470_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[20\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1197 net1198 vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__buf_2
X_14986_ net1121 vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09503__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_746 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16725_ clknet_leaf_173_wb_clk_i _02355_ _00421_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13937_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[4\] team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11310__B1 _07118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13552__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13868_ net1570 net983 _03770_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[5\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16656_ clknet_leaf_137_wb_clk_i _02286_ _00352_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12676__B net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15607_ net1169 vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__inv_2
X_12819_ net295 net2938 net486 vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__mux2_1
X_13799_ net1589 net974 net725 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[10\]
+ sky130_fd_sc_hd__and3_1
X_16587_ clknet_leaf_187_wb_clk_i _02217_ _00283_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08609__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18326_ net1317 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_56_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15538_ net1139 vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15469_ net1164 vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__inv_2
X_18257_ clknet_leaf_39_wb_clk_i _03486_ _01952_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_97_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17208_ clknet_leaf_29_wb_clk_i _02838_ _00904_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18188_ clknet_leaf_41_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[9\]
+ _01883_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09034__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold603 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net2017 sky130_fd_sc_hd__dlygate4sd3_1
Xhold614 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2028 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08242__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17139_ clknet_leaf_165_wb_clk_i _02769_ _00835_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold625 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net2039 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold636 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net2050 sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 net2061 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14315__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold658 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 net2072 sky130_fd_sc_hd__dlygate4sd3_1
X_09961_ _05895_ _05901_ _05988_ vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__or3_1
Xhold669 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2083 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08912_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[16\]
+ net648 net594 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[16\]
+ _04975_ vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12631__S _03682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09892_ _04428_ _05920_ vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__xnor2_4
X_08843_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[18\]
+ net814 net741 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__a22o_1
Xhold1303 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2717 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10352__A1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1314 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 net2728 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1325 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net2739 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1336 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net2750 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12629__A0 _03645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10004__X _06033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08774_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[19\]
+ net710 net649 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__a22o_1
Xhold1347 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 net2761 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1358 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 net2772 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1369 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net2783 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11301__B1 _07108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08848__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout456_A _03712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13462__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1198_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_74_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout623_A net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09326_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[8\]
+ net593 _05367_ _05373_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[8\]
+ sky130_fd_sc_hd__o22a_4
XFILLER_0_164_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12801__A0 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_153_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11604__B2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[21\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09273__A2 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09257_ net954 _04351_ _04269_ vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12806__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08481__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout411_X net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1153_X net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08208_ _04232_ net962 _04271_ _04156_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_170_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09188_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[10\]
+ net707 net632 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09025__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08139_ net1617 _04221_ _04225_ vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_79_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14306__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11150_ _07080_ _07114_ vssd1 vssd1 vccd1 vccd1 _07116_ sky130_fd_sc_hd__nor2_4
XANTENNA_fanout780_X net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13637__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10101_ _05350_ net361 vssd1 vssd1 vccd1 vccd1 _06129_ sky130_fd_sc_hd__or2_1
X_11081_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[4\] team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[3\]
+ vssd1 vssd1 vccd1 vccd1 _07048_ sky130_fd_sc_hd__nand2_1
XANTENNA__12541__S net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10032_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[13\] _04158_
+ _05923_ vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__or3_1
XANTENNA__09733__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14840_ net1201 vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_125_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14771_ net1213 vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__inv_2
XANTENNA_input17_A DAT_I[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11983_ _07719_ _07748_ vssd1 vssd1 vccd1 vccd1 _07795_ sky130_fd_sc_hd__or2_1
XANTENNA__08839__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13372__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13722_ net905 _06369_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[22\]
+ sky130_fd_sc_hd__and2_1
X_16510_ clknet_leaf_162_wb_clk_i _02140_ _00206_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10934_ net1043 _06343_ vssd1 vssd1 vccd1 vccd1 _06924_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17490_ clknet_leaf_36_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[25\]
+ _01186_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13653_ net2057 net331 net390 vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__mux2_1
X_16441_ clknet_leaf_9_wb_clk_i _02071_ _00137_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10865_ _06814_ _06861_ _06815_ vssd1 vssd1 vccd1 vccd1 _06862_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12604_ _03666_ net1746 net203 vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__mux2_1
X_16372_ clknet_leaf_111_wb_clk_i _02002_ _00068_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13584_ net2028 net304 net398 vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__mux2_1
X_10796_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[22\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06793_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09264__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18111_ clknet_leaf_55_wb_clk_i _03434_ _01807_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[28\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_143_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15323_ net1099 vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__inv_2
X_12535_ net1664 _03666_ net209 vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12716__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18042_ clknet_leaf_96_wb_clk_i _03380_ _01738_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_124_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15254_ net1096 vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__inv_2
X_12466_ net1629 _03666_ net212 vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__mux2_1
X_14205_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[9\] _04006_
+ vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11417_ net2970 _07323_ net1910 vssd1 vssd1 vccd1 vccd1 _07338_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15185_ net1188 vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12397_ net1674 _03666_ net217 vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08214__B net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14136_ net2306 net503 net911 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[19\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__09972__B1 _05924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11348_ net979 net508 net359 team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__a22o_1
X_18297__1389 vssd1 vssd1 vccd1 vccd1 net1389 _18297__1389/LO sky130_fd_sc_hd__conb_1
XANTENNA__13547__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14067_ _03934_ net979 team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__mux2_1
XANTENNA__12451__S net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11279_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[26\] _07119_
+ _07121_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[82\] _07239_
+ vssd1 vssd1 vccd1 vccd1 _07240_ sky130_fd_sc_hd__a221o_1
X_13018_ net300 net2225 net462 vssd1 vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17826_ clknet_leaf_92_wb_clk_i _03169_ _01522_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[72\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17757_ clknet_leaf_91_wb_clk_i _03100_ _01453_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_14969_ net1053 vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__inv_2
XANTENNA__09488__C1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13282__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16708_ clknet_leaf_179_wb_clk_i _02338_ _00404_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08490_ _04561_ _04563_ _04565_ _04567_ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__or4_2
XFILLER_0_77_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17688_ clknet_leaf_92_wb_clk_i _03031_ _01384_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[126\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08229__X _04312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13036__A0 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16639_ clknet_leaf_155_wb_clk_i _02269_ _00335_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_146_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09996__A _05034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10000__A _05165_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17986__Q net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11598__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09111_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[12\]
+ net777 net768 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18309_ net1401 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
XFILLER_0_115_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12626__S net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11530__S _07345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10270__B1 _04265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09042_ _05100_ vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09007__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold400 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[126\] vssd1 vssd1
+ vccd1 vccd1 net1814 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_192_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_192_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold411 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[97\] vssd1 vssd1
+ vccd1 vccd1 net1825 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout204_A _03681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold422 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[97\] vssd1 vssd1
+ vccd1 vccd1 net1836 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08899__X team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[17\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold433 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[48\] vssd1 vssd1
+ vccd1 vccd1 net1847 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[59\] vssd1 vssd1
+ vccd1 vccd1 net1858 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08766__B2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_121_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_121_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold455 net115 vssd1 vssd1 vccd1 vccd1 net1869 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold466 _03298_ vssd1 vssd1 vccd1 vccd1 net1880 sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[10\] vssd1
+ vssd1 vccd1 vccd1 net1891 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13457__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold488 net83 vssd1 vssd1 vccd1 vccd1 net1902 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout902 _04235_ vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__buf_2
X_09944_ _05933_ _05971_ _04925_ vssd1 vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__a21o_1
Xfanout913 net914 vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__buf_2
Xhold499 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[67\] vssd1 vssd1
+ vccd1 vccd1 net1913 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout924 net925 vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__clkbuf_2
Xfanout935 net937 vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__buf_2
Xfanout946 net949 vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__clkbuf_2
Xfanout957 net958 vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__clkbuf_2
X_09875_ _04677_ _05903_ vssd1 vssd1 vccd1 vccd1 _05904_ sky130_fd_sc_hd__nand2_1
XANTENNA_input9_A DAT_I[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout968 _04238_ vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__clkbuf_4
Xhold1100 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2514 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout979 team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[9\] vssd1 vssd1
+ vccd1 vccd1 net979 sky130_fd_sc_hd__buf_2
Xhold1111 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2525 sky130_fd_sc_hd__dlygate4sd3_1
X_18316__1408 vssd1 vssd1 vccd1 vccd1 net1408 _18316__1408/LO sky130_fd_sc_hd__conb_1
X_08826_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[18\]
+ net703 net682 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[18\]
+ _04894_ vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__a221o_1
Xhold1122 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net2536 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1133 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 net2547 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1144 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1155 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net2569 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1166 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2580 sky130_fd_sc_hd__dlygate4sd3_1
X_08757_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[21\]
+ net811 net739 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[21\]
+ _04828_ vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__a221o_1
Xhold1177 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1188 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net2602 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout740_A _04421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1199 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2613 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13192__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout838_A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout459_X net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08688_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[22\]
+ net712 net698 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__a22o_1
XANTENNA__09494__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18284__A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout626_X net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13578__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10650_ _06651_ _06654_ _04264_ vssd1 vssd1 vccd1 vccd1 _06655_ sky130_fd_sc_hd__a21oi_4
XANTENNA__09246__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09309_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[8\]
+ net848 net817 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__a22o_1
XANTENNA__12536__S _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10581_ _05817_ _05957_ _05285_ vssd1 vssd1 vccd1 vccd1 _06589_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12320_ _03611_ _03613_ _03608_ vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10261__B1 _06284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_39_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12251_ _08021_ _03514_ vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__and2b_1
XFILLER_0_121_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11202_ _07161_ _07163_ _07164_ _07166_ vssd1 vssd1 vccd1 vccd1 _07167_ sky130_fd_sc_hd__or4_1
XFILLER_0_82_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12182_ _07991_ _07992_ vssd1 vssd1 vccd1 vccd1 _07994_ sky130_fd_sc_hd__nor2_1
XANTENNA__13367__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11133_ _07072_ _07098_ vssd1 vssd1 vccd1 vccd1 _07099_ sky130_fd_sc_hd__nor2_4
X_16990_ clknet_leaf_162_wb_clk_i _02620_ _00686_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11064_ _07025_ _07029_ vssd1 vssd1 vccd1 vccd1 _07031_ sky130_fd_sc_hd__nand2_4
X_15941_ net1288 vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__inv_2
XANTENNA__09182__A1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ net364 net360 vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__nand2_1
X_15872_ net1264 vssd1 vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__inv_2
X_17611_ clknet_leaf_62_wb_clk_i _02982_ _01307_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_48_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14823_ net1176 vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__inv_2
XANTENNA_output123_A net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17542_ clknet_leaf_61_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[13\]
+ _01238_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11966_ _07741_ _07744_ _07742_ vssd1 vssd1 vccd1 vccd1 _07778_ sky130_fd_sc_hd__a21o_1
X_14754_ net1204 vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__inv_2
XANTENNA__10298__Y _06320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09485__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10739__B net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10917_ _06268_ _06909_ net1044 vssd1 vssd1 vccd1 vccd1 _06910_ sky130_fd_sc_hd__mux2_1
X_13705_ net900 _06672_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[5\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17473_ clknet_leaf_40_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[8\]
+ _01169_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11292__A2 _07100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14685_ net1092 vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__inv_2
XANTENNA__08693__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11897_ _07707_ _07708_ vssd1 vssd1 vccd1 vccd1 _07709_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08209__B net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16424_ clknet_leaf_197_wb_clk_i _02054_ _00120_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13636_ net2033 net248 net390 vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__mux2_1
X_10848_ _06842_ _06843_ _06837_ vssd1 vssd1 vccd1 vccd1 _06845_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_27_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09237__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12446__S _03670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16355_ clknet_leaf_192_wb_clk_i _01985_ _00051_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13567_ net2127 net237 net398 vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__mux2_1
XANTENNA__08445__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10779_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[30\] net1041 vssd1
+ vssd1 vccd1 vccd1 _06776_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_57_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12518_ net1932 _03646_ _03676_ vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__mux2_1
X_15306_ net1110 vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__inv_2
X_16286_ net1253 vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13498_ net2148 net222 net405 vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18025_ clknet_leaf_97_wb_clk_i _03364_ _01721_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12449_ net1724 _03646_ _03671_ vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__mux2_1
X_15237_ net1194 vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15168_ net1196 vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__inv_2
XANTENNA__13277__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14119_ _03950_ _03972_ _03982_ vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_1_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout209 _03676_ vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__buf_4
X_15099_ net1099 vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_66_Left_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09660_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[1\]
+ net787 _05671_ _05672_ _05678_ vssd1 vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__a2111oi_1
XTAP_TAPCELL_ROW_2_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08920__A1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08611_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[24\]
+ net649 net630 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[24\]
+ _04685_ vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__a221o_1
X_17809_ clknet_leaf_100_wb_clk_i _03152_ _01505_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09591_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[2\]
+ net760 _05602_ _05612_ _05616_ vssd1 vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_55_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08542_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[26\]
+ net843 net770 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_32_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_77_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09476__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12480__A1 _07789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08473_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[28\]
+ net593 _04542_ _04551_ vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_106_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_75_Left_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08436__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1063_A net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout419_A _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09025_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[14\]
+ net831 net791 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout207_X net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1230_A net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold230 net124 vssd1 vssd1 vccd1 vccd1 net1644 sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[115\] vssd1 vssd1
+ vccd1 vccd1 net1655 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold252 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[96\] vssd1 vssd1
+ vccd1 vccd1 net1666 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold263 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[90\] vssd1 vssd1
+ vccd1 vccd1 net1677 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout788_A _04400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13187__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold274 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[46\] vssd1 vssd1
+ vccd1 vccd1 net1688 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold285 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[34\] vssd1 vssd1
+ vccd1 vccd1 net1699 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold296 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[77\] vssd1 vssd1
+ vccd1 vccd1 net1710 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout710 _04290_ vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__clkbuf_8
Xfanout721 _04285_ vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__buf_6
Xfanout732 _07030_ vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_165_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09927_ _05378_ _05955_ _05939_ vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_leaf_71_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout743 net744 vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__buf_4
Xfanout754 net755 vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__clkbuf_4
Xfanout765 net767 vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08301__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout776 net777 vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__clkbuf_4
X_09858_ _05886_ vssd1 vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__inv_2
Xfanout787 _04400_ vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout798 net801 vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__buf_6
X_08809_ net571 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[19\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[19\] vssd1 vssd1 vccd1
+ vccd1 _04878_ sky130_fd_sc_hd__a21o_1
X_09789_ _05819_ vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout743_X net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11435__S net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11820_ _07630_ _07631_ vssd1 vssd1 vccd1 vccd1 _07632_ sky130_fd_sc_hd__nor2_1
X_11751_ net550 _07552_ _07558_ _07551_ vssd1 vssd1 vccd1 vccd1 _07563_ sky130_fd_sc_hd__a31o_1
XANTENNA__11274__A2 _07099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12471__A1 _03641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08675__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18296__1388 vssd1 vssd1 vccd1 vccd1 net1388 _18296__1388/LO sky130_fd_sc_hd__conb_1
XFILLER_0_95_354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13650__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10702_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[4\] net906 net897
+ _06703_ vssd1 vssd1 vccd1 vccd1 _06704_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_55_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14470_ net1231 vssd1 vssd1 vccd1 vccd1 _00100_ sky130_fd_sc_hd__inv_2
X_11682_ net70 net69 net41 net40 vssd1 vssd1 vccd1 vccd1 _07496_ sky130_fd_sc_hd__or4_1
XFILLER_0_138_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09219__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13421_ net1993 net313 net419 vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10633_ net2511 net294 net541 vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__mux2_1
XANTENNA__08427__B1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16140_ net1274 vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13352_ net295 net2533 net427 vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__mux2_1
X_10564_ _05826_ _05959_ vssd1 vssd1 vccd1 vccd1 _06573_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08045__A team_05_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10294__B _06316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12303_ _03569_ _03594_ _03597_ vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16071_ net1260 vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13283_ net293 net2517 net432 vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__mux2_1
X_10495_ _06061_ _05531_ vssd1 vssd1 vccd1 vccd1 _06508_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_20_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15022_ net1191 vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__inv_2
X_12234_ net354 _03510_ vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13097__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18250__Q team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12165_ _07927_ _07929_ _07971_ _07974_ _07976_ vssd1 vssd1 vccd1 vccd1 _07977_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_9_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11116_ _07073_ _07078_ vssd1 vssd1 vccd1 vccd1 _07083_ sky130_fd_sc_hd__nand2_2
X_16973_ clknet_leaf_160_wb_clk_i _02603_ _00669_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_12096_ _07864_ _07907_ vssd1 vssd1 vccd1 vccd1 _07908_ sky130_fd_sc_hd__nor2_1
X_15924_ net1293 vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__inv_2
X_11047_ _06846_ _07015_ net1044 vssd1 vssd1 vccd1 vccd1 _07016_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_30_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08363__C1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 DAT_I[16] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
X_15855_ net1294 vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14806_ net1091 vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15786_ net1295 vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__inv_2
X_12998_ net189 net2265 net461 vssd1 vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17525_ clknet_leaf_113_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[28\]
+ _01221_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12462__A1 _07798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14737_ net1189 vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__inv_2
XANTENNA__08666__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11949_ _07756_ _07757_ _07760_ vssd1 vssd1 vccd1 vccd1 _07761_ sky130_fd_sc_hd__a21o_1
XANTENNA__13560__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_116_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17456_ clknet_leaf_61_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[24\]
+ _01152_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14668_ net1071 vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12684__B net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16407_ clknet_leaf_143_wb_clk_i _02037_ _00103_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08418__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13619_ net2868 net315 net395 vssd1 vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__mux2_1
X_17387_ clknet_leaf_50_wb_clk_i net1429 _01083_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_14599_ net1104 vssd1 vssd1 vccd1 vccd1 _00229_ sky130_fd_sc_hd__inv_2
XANTENNA__10225__B1 _05924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11568__A3 _07422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16338_ net1119 vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18315__1407 vssd1 vssd1 vccd1 vccd1 net1407 _18315__1407/LO sky130_fd_sc_hd__conb_1
XANTENNA__09091__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16269_ net1115 vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__inv_2
XANTENNA__12904__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18008_ clknet_leaf_64_wb_clk_i _03347_ _01704_ vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire377_X net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09712_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[0\]
+ net950 net1014 net929 vssd1 vssd1 vccd1 vccd1 _05744_ sky130_fd_sc_hd__and4_1
X_09643_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[1\]
+ net942 net938 _04418_ vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__and4_1
XANTENNA_clkbuf_leaf_155_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10700__A1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout369_A _05577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09574_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[2\]
+ net941 net1013 net927 vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__and4_1
XFILLER_0_136_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09449__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08525_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[26\]
+ net714 net600 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[26\]
+ _04601_ vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__a221o_1
XANTENNA__11256__A2 _07092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout536_A net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13470__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1278_A net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08456_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[28\]
+ net831 net800 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[28\]
+ _04534_ vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__a221o_1
XFILLER_0_129_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08387_ net380 _04466_ vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout703_A _04292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10216__B1 _06237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09082__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09621__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12814__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09008_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[14\]
+ net619 net615 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[14\]
+ _05068_ vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_167_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10280_ _05903_ _06051_ _06302_ _06056_ _05905_ vssd1 vssd1 vccd1 vccd1 _06303_ sky130_fd_sc_hd__a32o_1
XANTENNA__08152__X _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10519__A1 _06049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout693_X net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14314__B team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[20\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_194_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08312__B net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout860_X net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout958_X net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout540 net541 vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__clkbuf_8
Xfanout551 net553 vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13645__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout562 _03692_ vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__clkbuf_2
X_13970_ _03840_ _03841_ _03821_ vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__o21a_1
Xfanout573 _04343_ vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14330__A team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09688__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout595 net597 vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__clkbuf_8
X_12921_ net314 net2442 net475 vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__mux2_1
XANTENNA__08896__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08360__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15640_ net1246 vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__inv_2
X_12852_ net294 net2330 net482 vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11803_ _07607_ _07609_ _07611_ _07612_ _07613_ vssd1 vssd1 vccd1 vccd1 _07615_ sky130_fd_sc_hd__a32o_2
XANTENNA__11247__A2 _07102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12444__A1 _03651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12783_ net298 net2598 net490 vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__mux2_1
XANTENNA__08648__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15571_ net1282 vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__inv_2
XANTENNA__13380__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17310_ clknet_leaf_178_wb_clk_i _02940_ _01006_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_2
X_11734_ _07542_ _07543_ _07544_ vssd1 vssd1 vccd1 vccd1 _07546_ sky130_fd_sc_hd__nor3_1
X_14522_ net1058 vssd1 vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18290_ net1382 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
XFILLER_0_68_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09860__A2 _05881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17241_ clknet_leaf_9_wb_clk_i _02871_ _00937_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11665_ net28 net990 net917 net1865 vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_25_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14453_ net1060 vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10207__B1 _06055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10616_ _05378_ _05955_ vssd1 vssd1 vccd1 vccd1 _06622_ sky130_fd_sc_hd__xnor2_1
X_13404_ net2580 net227 net418 vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__mux2_1
X_14384_ net1504 vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09073__B1 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17172_ clknet_leaf_120_wb_clk_i _02802_ _00868_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11596_ net128 net1011 net346 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16123_ net1136 vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__inv_2
X_13335_ net238 net2620 net426 vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__mux2_1
X_10547_ _05189_ _05828_ vssd1 vssd1 vccd1 vccd1 _06557_ sky130_fd_sc_hd__xor2_2
XFILLER_0_122_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08820__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12724__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09158__X _05213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16054_ net1262 vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__inv_2
X_13266_ net218 net2287 net434 vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__mux2_1
X_10478_ _06338_ _06491_ net370 vssd1 vssd1 vccd1 vccd1 _06492_ sky130_fd_sc_hd__mux2_1
X_12217_ _08022_ _03510_ vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__nand2_4
X_15005_ net1090 vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13197_ _06247_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[28\]
+ net352 vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__mux2_1
XANTENNA__08222__B net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12148_ _07950_ _07958_ _07911_ vssd1 vssd1 vccd1 vccd1 _07960_ sky130_fd_sc_hd__a21boi_2
XANTENNA__10391__C1 _05924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13555__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12079_ _07888_ _07890_ vssd1 vssd1 vccd1 vccd1 _07891_ sky130_fd_sc_hd__and2_1
X_16956_ clknet_leaf_154_wb_clk_i _02586_ _00652_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08336__C1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[22\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12679__B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15907_ net1301 vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_139_Right_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16887_ clknet_leaf_146_wb_clk_i _02517_ _00583_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08887__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08351__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15838_ net1273 vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12435__A1 _07836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11238__A2 _07102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08639__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15769_ net1276 vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13290__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08310_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[31\]
+ net811 net807 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[31\]
+ _04389_ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_47_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17508_ clknet_leaf_114_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[11\]
+ _01204_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_09290_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[8\]
+ net685 net635 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[8\]
+ _05332_ vssd1 vssd1 vccd1 vccd1 _05339_ sky130_fd_sc_hd__a221o_1
XANTENNA__08237__X _04320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08241_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[31\]
+ net688 net657 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17439_ clknet_leaf_65_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[7\]
+ _01135_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08172_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[9\] _04249_
+ vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_95_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12634__S _03682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_99_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_132_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__buf_2
Xoutput121 net121 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__buf_2
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput132 net132 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__buf_2
Xoutput143 net143 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_28_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xoutput154 net154 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__clkbuf_4
Xoutput165 net165 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_110_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1026_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18295__1387 vssd1 vssd1 vccd1 vccd1 net1387 _18295__1387/LO sky130_fd_sc_hd__conb_1
XFILLER_0_100_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput176 net176 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__clkbuf_4
Xoutput187 net187 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13465__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout486_A _03703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08590__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10134__C1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout653_A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09626_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[2\]
+ net665 _05637_ _05648_ _05651_ vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_108_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11229__A2 _07092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09557_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[3\]
+ net629 _05593_ net719 vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout441_X net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout820_A net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12809__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09827__C1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout539_X net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08508_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[27\]
+ net772 net761 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[27\]
+ _04585_ vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__a221o_1
X_09488_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[4\]
+ net799 _05527_ net855 vssd1 vssd1 vccd1 vccd1 _05528_ sky130_fd_sc_hd__a211o_1
XFILLER_0_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09842__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08439_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[28\]
+ net705 net654 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_156_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout706_X net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11450_ _07346_ _07359_ _07358_ vssd1 vssd1 vccd1 vccd1 _07361_ sky130_fd_sc_hd__o21a_1
XANTENNA__10417__A2_N _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09055__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10401_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[20\] _06096_ vssd1
+ vssd1 vccd1 vccd1 _06419_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11381_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[6\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[5\]
+ vssd1 vssd1 vccd1 vccd1 _07312_ sky130_fd_sc_hd__nand2_1
XANTENNA__08802__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Left_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13120_ net318 net2190 net448 vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__mux2_1
X_10332_ _06032_ net338 net333 _06047_ vssd1 vssd1 vccd1 vccd1 _06353_ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13051_ net301 net2358 net459 vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__mux2_1
X_10263_ _06155_ _06170_ net531 vssd1 vssd1 vccd1 vccd1 _06287_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12002_ _07477_ _07517_ _07800_ _07813_ _07796_ vssd1 vssd1 vccd1 vccd1 _07814_ sky130_fd_sc_hd__a221o_1
Xfanout1302 net1303 vssd1 vssd1 vccd1 vccd1 net1302 sky130_fd_sc_hd__buf_4
XANTENNA_input47_A wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10194_ net893 _06219_ vssd1 vssd1 vccd1 vccd1 _06220_ sky130_fd_sc_hd__nor2_1
Xfanout1313 net38 vssd1 vssd1 vccd1 vccd1 net1313 sky130_fd_sc_hd__buf_6
XANTENNA__13375__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16810_ clknet_leaf_17_wb_clk_i _02440_ _00506_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08581__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17790_ clknet_leaf_84_wb_clk_i _03133_ _01486_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[100\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout370 net372 vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__buf_4
X_16741_ clknet_leaf_22_wb_clk_i _02371_ _00437_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout392 _03732_ vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__buf_6
X_13953_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[9\] _03825_ vssd1
+ vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__xor2_1
XANTENNA__08869__B1 _04318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18314__1406 vssd1 vssd1 vccd1 vccd1 net1406 _18314__1406/LO sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_21_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12904_ net227 net2827 net475 vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__mux2_1
X_16672_ clknet_leaf_132_wb_clk_i _02302_ _00368_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13884_ net1579 net982 _03778_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[13\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18411_ net915 vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__clkbuf_1
X_15623_ net1160 vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12835_ net240 net2495 net482 vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12719__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10428__B1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18342_ net1331 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
X_15554_ net1123 vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12766_ net245 net2293 net491 vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__mux2_1
XANTENNA__09294__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09833__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14505_ net1214 vssd1 vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__inv_2
X_18273_ clknet_leaf_36_wb_clk_i _03502_ _01968_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[27\]
+ sky130_fd_sc_hd__dfrtp_4
X_11717_ net356 _07527_ vssd1 vssd1 vccd1 vccd1 _07529_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15485_ net1147 vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__inv_2
X_12697_ net225 net2597 net497 vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__mux2_1
XANTENNA__08217__B net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17224_ clknet_leaf_196_wb_clk_i _02854_ _00920_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11648_ net15 net991 net918 net1942 vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__a22o_1
X_14436_ net1226 vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__inv_2
XANTENNA__09046__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput12 DAT_I[19] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
Xinput23 DAT_I[29] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
Xinput34 gpio_in[34] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_1
Xinput45 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17155_ clknet_leaf_199_wb_clk_i _02785_ _00851_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11579_ net1935 net1005 _07398_ net357 vssd1 vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__a22o_1
XANTENNA__12454__S net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14367_ _04094_ _04138_ _04139_ vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__or3_1
Xinput56 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput67 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__clkbuf_1
Xhold807 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net2221 sky130_fd_sc_hd__dlygate4sd3_1
X_16106_ net1310 vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__inv_2
XANTENNA__10600__B1 _04279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13318_ net2068 net300 net429 vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__mux2_1
Xhold818 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2232 sky130_fd_sc_hd__dlygate4sd3_1
Xhold829 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2243 sky130_fd_sc_hd__dlygate4sd3_1
X_17086_ clknet_leaf_163_wb_clk_i _02716_ _00782_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_14298_ net379 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16037_ net1250 vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__inv_2
X_13249_ net281 net2241 net437 vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13285__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08572__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1507 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2921 sky130_fd_sc_hd__dlygate4sd3_1
X_08790_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[19\]
+ net777 net768 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__a22o_1
X_17988_ clknet_leaf_83_wb_clk_i _03327_ _01684_ vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__dfrtp_1
Xhold1518 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 net2932 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1529 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net2943 sky130_fd_sc_hd__dlygate4sd3_1
X_16939_ clknet_leaf_187_wb_clk_i _02569_ _00635_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12656__A1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[11\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10667__B1 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_146_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_146_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09999__A _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09411_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[6\]
+ net841 net818 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[6\]
+ _05454_ vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12629__S net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10938__A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09342_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[7\]
+ net688 net657 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[7\]
+ _05388_ vssd1 vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_138_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09285__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09824__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09273_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[9\]
+ net838 net779 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[9\]
+ _05322_ vssd1 vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_62_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout234_A net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11550__A_N _07396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08224_ net879 net872 net865 vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__and3_1
XFILLER_0_145_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08155_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[2\] _04229_
+ _04236_ vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__and3_1
XANTENNA__10673__A _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout401_A net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14145__A team_05_WB.instance_to_wrap.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12592__A0 _03614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1143_A net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08086_ net1025 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[18\]
+ net971 _04192_ vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1310_A net1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout391_X net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13195__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout489_X net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout868_A _04289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08563__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08988_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[15\]
+ net845 net771 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout656_X net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08315__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10950_ net1042 _06401_ vssd1 vssd1 vccd1 vccd1 _06937_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_127_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09609_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[2\]
+ net886 net875 net870 vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_158_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10881_ _06789_ _06877_ _06788_ vssd1 vssd1 vccd1 vccd1 _06878_ sky130_fd_sc_hd__a21boi_1
XANTENNA_fanout823_X net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12539__S _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12620_ net1679 _07793_ _03682_ vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09276__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09815__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12551_ _03657_ net1784 net205 vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11502_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[19\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[19\]
+ net1031 vssd1 vssd1 vccd1 vccd1 _07413_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12482_ net1820 _03657_ net211 vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__mux2_1
X_15270_ net1209 vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__inv_2
XANTENNA__09028__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11433_ net1050 net1049 vssd1 vssd1 vccd1 vccd1 _07346_ sky130_fd_sc_hd__or2_4
X_14221_ team_05_WB.instance_to_wrap.total_design.keypad0.counter\[0\] team_05_WB.instance_to_wrap.total_design.keypad0.counter\[1\]
+ team_05_WB.instance_to_wrap.total_design.keypad0.counter\[2\] vssd1 vssd1 vccd1
+ vccd1 _04017_ sky130_fd_sc_hd__and3_1
XFILLER_0_151_524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10189__A2 _06214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14152_ _03809_ _03994_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[1\]
+ sky130_fd_sc_hd__nor2_1
X_11364_ _07286_ _07291_ _07292_ _07302_ vssd1 vssd1 vccd1 vccd1 _07304_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_81_1036 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13103_ net232 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[23\]
+ net450 vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__mux2_1
XANTENNA__14324__A1 _05442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10315_ _05634_ _06336_ _06334_ vssd1 vssd1 vccd1 vccd1 _06337_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_104_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14083_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[10\] net980 _03801_
+ vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__o21ai_2
XANTENNA__14324__B2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[5\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11295_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[25\] _07119_
+ _07120_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[33\] vssd1 vssd1
+ vccd1 vccd1 _07255_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17911_ clknet_leaf_88_wb_clk_i _03254_ _01607_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13034_ net242 net2768 net458 vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__mux2_1
X_10246_ net383 _06270_ vssd1 vssd1 vccd1 vccd1 _06271_ sky130_fd_sc_hd__and2_1
XANTENNA__09200__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1110 net1111 vssd1 vssd1 vccd1 vccd1 net1110 sky130_fd_sc_hd__clkbuf_4
Xfanout1121 net1127 vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__buf_4
X_17842_ clknet_leaf_91_wb_clk_i _03185_ _01538_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[88\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1132 net1133 vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__clkbuf_4
X_10177_ _06073_ _06192_ _06203_ vssd1 vssd1 vccd1 vccd1 _06204_ sky130_fd_sc_hd__o21a_1
Xfanout1143 net1151 vssd1 vssd1 vccd1 vccd1 net1143 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1081 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1154 net1162 vssd1 vssd1 vccd1 vccd1 net1154 sky130_fd_sc_hd__buf_4
Xfanout1165 net1175 vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__clkbuf_4
Xfanout1176 net1177 vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__buf_4
X_17773_ clknet_leaf_102_wb_clk_i _03116_ _01469_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1187 net1190 vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__buf_4
X_14985_ net1221 vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__inv_2
Xfanout1198 net1211 vssd1 vssd1 vccd1 vccd1 net1198 sky130_fd_sc_hd__buf_2
XANTENNA__10649__B1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16724_ clknet_leaf_119_wb_clk_i _02354_ _00420_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_13936_ _03805_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[2\] vssd1
+ vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__and2b_1
XFILLER_0_89_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16655_ clknet_leaf_136_wb_clk_i _02285_ _00351_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13867_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[5\]
+ net559 net575 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[5\]
+ net986 vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__a221o_1
XANTENNA__12449__S _03671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15606_ net1258 vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_83_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12818_ net299 net2544 net487 vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__mux2_1
XANTENNA__09267__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16586_ clknet_leaf_195_wb_clk_i _02216_ _00282_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_146_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13798_ net1415 net974 net725 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[9\]
+ sky130_fd_sc_hd__and3_1
X_18325_ net1316 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
X_18294__1386 vssd1 vssd1 vccd1 vccd1 net1386 _18294__1386/LO sky130_fd_sc_hd__conb_1
X_15537_ net1140 vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12749_ net286 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[10\]
+ net492 vssd1 vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10196__C _05801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18256_ clknet_leaf_41_wb_clk_i _03485_ _01951_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_13_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13788__B _03748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15468_ net1164 vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17207_ clknet_leaf_145_wb_clk_i _02837_ _00903_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14419_ net1213 vssd1 vssd1 vccd1 vccd1 _00049_ sky130_fd_sc_hd__inv_2
XFILLER_0_163_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18187_ clknet_leaf_40_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[8\]
+ _01882_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15399_ net1242 vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__inv_2
X_17138_ clknet_leaf_125_wb_clk_i _02768_ _00834_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold604 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2018 sky130_fd_sc_hd__dlygate4sd3_1
Xhold615 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2029 sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2040 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold637 net103 vssd1 vssd1 vccd1 vccd1 net2051 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14315__A1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08793__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold648 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2062 sky130_fd_sc_hd__dlygate4sd3_1
X_09960_ _05895_ _05988_ vssd1 vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__nor2_1
Xhold659 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2073 sky130_fd_sc_hd__dlygate4sd3_1
X_17069_ clknet_leaf_160_wb_clk_i _02699_ _00765_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14315__B2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[18\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12912__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16180__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08911_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[16\]
+ net711 net682 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__a22o_1
X_09891_ _04470_ _05919_ _04468_ vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08545__A2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08842_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[18\]
+ net845 net829 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[18\]
+ _04909_ vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__a221o_1
Xhold1304 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1315 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net2729 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1326 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2740 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08773_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[19\]
+ net625 net606 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[19\]
+ _04843_ vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__a221o_1
Xhold1337 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2751 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1348 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2762 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1359 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2773 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15524__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout351_A _03717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1093_A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout449_A _03714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10020__X _06049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09325_ _05368_ _05369_ _05370_ _05372_ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__or4_1
XANTENNA__11604__A2 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1260_A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout237_X net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout616_A _04318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09256_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[27\] _04350_
+ net953 vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08207_ net884 net870 net868 vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_43_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09187_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[10\]
+ net660 net625 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_170_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout404_X net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12565__A0 _03604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18313__1405 vssd1 vssd1 vccd1 vccd1 net1405 _18313__1405/LO sky130_fd_sc_hd__conb_1
X_08138_ _04216_ _04224_ _04218_ vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__a21o_1
XFILLER_0_133_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09430__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout985_A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08784__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14306__A1 _04656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08069_ net1024 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__and2b_1
XANTENNA__14306__B2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[24\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1313_X net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12822__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10591__A2 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10100_ _06126_ _06127_ vssd1 vssd1 vccd1 vccd1 _06128_ sky130_fd_sc_hd__nand2_1
X_11080_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[1\] team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[2\]
+ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[0\] vssd1 vssd1
+ vccd1 vccd1 _07047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout773_X net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14322__B team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[16\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08536__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10031_ net531 _06059_ vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__nand2_2
XFILLER_0_76_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout940_X net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11962__A team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13653__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14770_ net1235 vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__inv_2
X_11982_ _07789_ _07791_ _07793_ vssd1 vssd1 vccd1 vccd1 _07794_ sky130_fd_sc_hd__nand3_1
XANTENNA__09497__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13721_ _04235_ _06387_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[21\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10933_ _06790_ _06877_ vssd1 vssd1 vccd1 vccd1 _06923_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_169_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16440_ clknet_leaf_33_wb_clk_i _02070_ _00136_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10864_ _06816_ _06860_ vssd1 vssd1 vccd1 vccd1 _06861_ sky130_fd_sc_hd__or2_1
X_13652_ net2044 net314 net391 vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__mux2_1
XANTENNA__08048__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12603_ _03665_ net1832 _03681_ vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__mux2_1
X_16371_ clknet_leaf_165_wb_clk_i _02001_ _00067_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10795_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[23\] net1040 vssd1
+ vssd1 vccd1 vccd1 _06792_ sky130_fd_sc_hd__or2_1
X_13583_ net2106 net296 net399 vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__mux2_1
XANTENNA__12793__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[10\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18110_ clknet_leaf_55_wb_clk_i _03433_ _01806_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[27\]
+ sky130_fd_sc_hd__dfrtp_4
X_15322_ net1053 vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12534_ net1837 _03665_ net208 vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08335__X _04417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18041_ clknet_leaf_95_wb_clk_i _03379_ _01737_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__18253__Q team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15253_ net1079 vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__inv_2
X_12465_ net1728 _03665_ _03671_ vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__mux2_1
XANTENNA__12556__A0 _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08054__Y _04174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14204_ _04006_ net728 _04005_ vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__and3b_1
X_11416_ net1862 _07324_ vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__xor2_1
XFILLER_0_62_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12396_ _03531_ _03536_ _03540_ net354 _07914_ vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__a32o_2
X_15184_ net1092 vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__inv_2
XANTENNA__10567__C1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08214__C net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11347_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[10\] net508 net359
+ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[6\] vssd1 vssd1 vccd1
+ vccd1 _03393_ sky130_fd_sc_hd__a22o_1
X_14135_ team_05_WB.instance_to_wrap.CPU_DAT_O\[18\] net505 net912 vssd1 vssd1 vccd1
+ vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[18\] sky130_fd_sc_hd__and3_1
XANTENNA__09972__A1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08775__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12732__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11278_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[34\] _07120_
+ _07237_ _07238_ vssd1 vssd1 vccd1 vccd1 _07239_ sky130_fd_sc_hd__a211o_1
X_14066_ net979 net980 vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__nand2_1
XANTENNA__08527__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10229_ _06252_ _06253_ net371 vssd1 vssd1 vccd1 vccd1 _06254_ sky130_fd_sc_hd__mux2_1
X_13017_ net288 net2234 net460 vssd1 vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__mux2_1
XANTENNA__11531__A1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08230__B net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17825_ clknet_leaf_100_wb_clk_i _03168_ _01521_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[71\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_33_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[9\]
+ vssd1 vssd1 vccd1 vccd1 net1415 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_85_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13563__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17756_ clknet_leaf_83_wb_clk_i _03099_ _01452_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_22_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13790__C net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14968_ net1244 vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__inv_2
XANTENNA__12687__B net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11591__B _07452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16707_ clknet_leaf_198_wb_clk_i _02337_ _00403_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13919_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[31\]
+ net561 net577 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[31\]
+ net985 vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__a221o_1
XANTENNA__11295__B1 _07120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17687_ clknet_leaf_89_wb_clk_i _03030_ _01383_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[125\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14899_ net1212 vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_18_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16638_ clknet_leaf_184_wb_clk_i _02268_ _00334_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16569_ clknet_leaf_9_wb_clk_i _02199_ _00265_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16175__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12907__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11598__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09110_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[24\] net968
+ net954 _05166_ _04345_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[12\]
+ sky130_fd_sc_hd__a221o_1
X_18308_ net1400 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
XFILLER_0_44_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09041_ net571 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[14\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[14\] vssd1 vssd1 vccd1
+ vccd1 _05100_ sky130_fd_sc_hd__a21o_1
X_18239_ clknet_leaf_57_wb_clk_i net1512 _01934_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__18390__A net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12547__A0 _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold401 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[9\] vssd1 vssd1
+ vccd1 vccd1 net1815 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09412__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold412 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[86\] vssd1 vssd1
+ vccd1 vccd1 net1826 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[7\] vssd1 vssd1
+ vccd1 vccd1 net1837 sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[52\] vssd1 vssd1
+ vccd1 vccd1 net1848 sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[8\] vssd1 vssd1
+ vccd1 vccd1 net1859 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12642__S _03682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold456 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[2\] vssd1 vssd1
+ vccd1 vccd1 net1870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[18\] vssd1 vssd1
+ vccd1 vccd1 net1881 sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[48\] vssd1 vssd1
+ vccd1 vccd1 net1892 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold489 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[111\] vssd1 vssd1
+ vccd1 vccd1 net1903 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09943_ _05933_ _05971_ _04925_ vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_61_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout903 net904 vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__buf_4
Xfanout914 net915 vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17507__Q team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[10\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout925 net926 vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__buf_2
XANTENNA__08518__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_0_wb_clk_i_X clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout399_A _03731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout936 net937 vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__buf_2
X_09874_ _04656_ _04676_ vssd1 vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_161_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_161_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout947 net949 vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_146_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout958 net959 vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_146_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout969 net973 vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__buf_2
Xhold1101 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 net2515 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1106_A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1112 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[14\] vssd1 vssd1
+ vccd1 vccd1 net2526 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09191__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08825_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[18\]
+ net683 net648 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__a22o_1
Xhold1123 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1134 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2548 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13473__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1145 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2559 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1156 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2570 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1167 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2581 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09479__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08756_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[21\]
+ net842 net823 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__a22o_1
Xhold1178 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net2592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1189 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net2603 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout733_A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08687_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[22\]
+ net684 net634 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout900_A net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12817__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout619_X net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13061__X _03713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09308_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[8\]
+ net843 net835 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05356_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10580_ net2353 net293 net539 vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__mux2_1
XANTENNA__08155__X _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09239_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[9\]
+ net709 net642 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__a22o_1
XANTENNA__13221__B net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12250_ _08009_ _08020_ _03543_ _08019_ vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_118_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout890_X net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09403__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout988_X net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11201_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[102\] _07123_
+ _07165_ _07069_ vssd1 vssd1 vccd1 vccd1 _07166_ sky130_fd_sc_hd__a211o_1
XANTENNA__11210__B1 _07130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08757__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13648__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12181_ _07992_ vssd1 vssd1 vccd1 vccd1 _07993_ sky130_fd_sc_hd__inv_2
XANTENNA__12552__S _03678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14333__A _05768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11132_ _07059_ _07075_ vssd1 vssd1 vccd1 vccd1 _07098_ sky130_fd_sc_hd__nand2_2
Xhold990 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2404 sky130_fd_sc_hd__dlygate4sd3_1
X_11063_ _07025_ _07029_ vssd1 vssd1 vccd1 vccd1 _07030_ sky130_fd_sc_hd__and2_1
X_15940_ net1296 vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__inv_2
X_18293__1385 vssd1 vssd1 vccd1 vccd1 net1385 _18293__1385/LO sky130_fd_sc_hd__conb_1
X_10014_ _04818_ net367 vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__nand2_1
XANTENNA__09182__A2 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15871_ net1292 vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__inv_2
XANTENNA__08113__A_N net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17610_ clknet_leaf_61_wb_clk_i _02981_ _01306_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13383__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14822_ net1209 vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__inv_2
XANTENNA__10579__Y _06588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17541_ clknet_leaf_61_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[12\]
+ _01237_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11277__B1 _07115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14753_ net1236 vssd1 vssd1 vccd1 vccd1 _00383_ sky130_fd_sc_hd__inv_2
X_11965_ _07767_ _07769_ _07773_ _07776_ _07765_ vssd1 vssd1 vccd1 vccd1 _07777_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_99_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output116_A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08049__Y _04170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13704_ net901 _06691_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[4\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_80_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10916_ _06881_ _06908_ vssd1 vssd1 vccd1 vccd1 _06909_ sky130_fd_sc_hd__xnor2_1
X_17472_ clknet_leaf_40_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[7\]
+ _01168_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_106_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_6_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14684_ net1074 vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__inv_2
XANTENNA__10101__A _05350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11896_ _07672_ _07678_ vssd1 vssd1 vccd1 vccd1 _07708_ sky130_fd_sc_hd__xor2_2
X_16423_ clknet_leaf_201_wb_clk_i _02053_ _00119_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08209__C net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13635_ net2029 net228 net391 vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__mux2_1
XANTENNA__10595__X _06603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10847_ _06837_ _06842_ _06843_ vssd1 vssd1 vccd1 vccd1 _06844_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16354_ clknet_leaf_8_wb_clk_i _01984_ _00050_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13566_ net2327 net238 net399 vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__mux2_1
X_10778_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[30\] net1041 vssd1
+ vssd1 vccd1 vccd1 _06775_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_4_Left_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10252__A1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15305_ net1221 vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__inv_2
X_12517_ _07793_ net1905 _03675_ vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__mux2_1
X_16285_ net1254 vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__inv_2
XANTENNA__10247__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13497_ net2064 net220 net406 vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08225__B net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18024_ clknet_leaf_96_wb_clk_i _03363_ _01720_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_15236_ net1230 vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__inv_2
X_12448_ net1807 _07793_ _03670_ vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13558__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08748__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12462__S _03670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15167_ net1179 vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__inv_2
X_12379_ net1708 _03644_ net216 vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__mux2_1
XANTENNA__12315__X _03610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10555__A2 _06237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14118_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[15\] _04159_ _03868_
+ _03981_ vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15098_ net1056 vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__inv_2
X_14049_ _03915_ _03917_ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_145_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_4__f_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08381__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13293__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08920__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08610_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[24\]
+ net706 net613 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17808_ clknet_leaf_104_wb_clk_i _03151_ _01504_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[118\]
+ sky130_fd_sc_hd__dfrtp_1
X_09590_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[2\]
+ net748 _05604_ _05619_ _05621_ vssd1 vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11268__B1 _07128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17739_ clknet_leaf_89_wb_clk_i _03082_ _01435_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_141_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18312__1404 vssd1 vssd1 vccd1 vccd1 net1404 _18312__1404/LO sky130_fd_sc_hd__conb_1
X_08541_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[26\]
+ net792 net776 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__a22o_1
XANTENNA__12210__B net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08472_ _04544_ _04546_ _04548_ _04550_ vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__or4_1
XFILLER_0_148_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09800__A _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12637__S _03683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11440__B1 team_05_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08987__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10157__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout314_A net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1056_A net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09024_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[14\]
+ net820 net808 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[14\]
+ _05083_ vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13468__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold220 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[64\] vssd1 vssd1
+ vccd1 vccd1 net1634 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08739__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12372__S _07852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold231 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[107\] vssd1 vssd1
+ vccd1 vccd1 net1645 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold242 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[25\] vssd1 vssd1
+ vccd1 vccd1 net1656 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_184_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1223_A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold253 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[25\]
+ vssd1 vssd1 vccd1 vccd1 net1667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[29\] vssd1 vssd1
+ vccd1 vccd1 net1678 sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[78\] vssd1 vssd1
+ vccd1 vccd1 net1689 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08151__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold286 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[84\] vssd1 vssd1
+ vccd1 vccd1 net1700 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout683_A net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout700 _04293_ vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10951__C1 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold297 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[15\] vssd1 vssd1
+ vccd1 vccd1 net1711 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout711 _04288_ vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__buf_6
X_09926_ _05423_ _05954_ _05940_ vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__a21oi_2
Xfanout722 _04285_ vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_165_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1011_X net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout733 net736 vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__clkbuf_8
Xfanout744 _04419_ vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__buf_4
Xfanout755 _04414_ vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09164__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout766 net767 vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__clkbuf_4
X_09857_ _04839_ _05885_ vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__and2_4
Xfanout777 _04404_ vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__buf_4
XANTENNA_fanout850_A _04370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout788 _04400_ vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout471_X net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08372__B1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout799 net801 vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout948_A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08808_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[19\]
+ net590 _04874_ _04877_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[19\]
+ sky130_fd_sc_hd__o22a_4
XANTENNA__08911__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09788_ _05331_ _05818_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__nand2_1
XANTENNA__11259__B1 _07126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08739_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[21\]
+ net688 net595 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout736_X net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15712__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11750_ _07547_ _07561_ vssd1 vssd1 vccd1 vccd1 _07562_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10701_ _06086_ _06702_ vssd1 vssd1 vccd1 vccd1 _06703_ sky130_fd_sc_hd__or2_1
X_11681_ net50 net39 net64 net61 vssd1 vssd1 vccd1 vccd1 _07495_ sky130_fd_sc_hd__or4_1
XANTENNA__12547__S net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11451__S net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14328__A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13420_ net2319 net319 net418 vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__mux2_1
X_10632_ _04264_ _06637_ vssd1 vssd1 vccd1 vccd1 _06638_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08326__A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10563_ _05822_ _05827_ vssd1 vssd1 vccd1 vccd1 _06572_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_24_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08978__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13351_ net299 net2914 net426 vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12302_ _03569_ _03594_ _03511_ vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__o21ai_1
X_16070_ net1260 vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__inv_2
XFILLER_0_161_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10494_ _04157_ net1018 _05056_ vssd1 vssd1 vccd1 vccd1 _06507_ sky130_fd_sc_hd__mux2_1
X_13282_ net280 net2136 net433 vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13378__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15021_ net1087 vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__inv_2
X_12233_ _03520_ _03526_ _03523_ vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__a21o_1
XFILLER_0_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10537__A2 _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12164_ _07920_ _07962_ _07969_ vssd1 vssd1 vccd1 vccd1 _07976_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_9_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11115_ _07072_ _07081_ vssd1 vssd1 vccd1 vccd1 _07082_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_9_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16972_ clknet_leaf_0_wb_clk_i _02602_ _00668_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_12095_ _07895_ _07903_ vssd1 vssd1 vccd1 vccd1 _07907_ sky130_fd_sc_hd__xnor2_2
X_15923_ net1304 vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__inv_2
X_11046_ _06835_ _06836_ _06845_ vssd1 vssd1 vccd1 vccd1 _07015_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_30_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15854_ net1256 vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__inv_2
XANTENNA__09604__B net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14805_ net1060 vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__inv_2
X_15785_ net1265 vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__inv_2
X_12997_ net195 net2322 net462 vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17524_ clknet_leaf_113_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[27\]
+ _01220_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[27\]
+ sky130_fd_sc_hd__dfrtp_4
X_14736_ net1102 vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11948_ _07733_ _07759_ _07739_ vssd1 vssd1 vccd1 vccd1 _07760_ sky130_fd_sc_hd__o21a_1
XFILLER_0_146_5 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17455_ clknet_leaf_57_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[23\]
+ _01151_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10473__B2 _06355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12457__S _03671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14667_ net1067 vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__inv_2
X_11879_ net549 _07690_ vssd1 vssd1 vccd1 vccd1 _07691_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16406_ clknet_leaf_142_wb_clk_i _02036_ _00102_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13618_ net2071 net319 net394 vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__mux2_1
X_17386_ clknet_leaf_49_wb_clk_i net1418 _01082_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_14598_ net1230 vssd1 vssd1 vccd1 vccd1 _00228_ sky130_fd_sc_hd__inv_2
X_16337_ net1117 vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__inv_2
XANTENNA__08969__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13549_ net2759 net300 net402 vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16268_ net1129 vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__inv_2
XANTENNA__10772__Y _06769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08159__A_N team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18007_ clknet_leaf_64_wb_clk_i _03346_ _01703_ vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13288__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15219_ net1213 vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16199_ net1146 vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__inv_2
XANTENNA__12045__X _07857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09394__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12920__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10006__A net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09146__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09711_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[0\]
+ net1017 net944 net934 vssd1 vssd1 vccd1 vccd1 _05743_ sky130_fd_sc_hd__and4_1
XANTENNA__08354__B1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09642_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[1\]
+ net940 net1013 net924 vssd1 vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__and4_1
XANTENNA__10700__A2 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09573_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[2\]
+ net1015 net941 net924 vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__and4_1
XFILLER_0_77_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08524_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[26\]
+ net697 net678 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08455_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[28\]
+ net762 net753 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__a22o_1
XANTENNA__17520__Q team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[23\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08386_ net570 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[30\]
+ _04362_ vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18292__1384 vssd1 vssd1 vccd1 vccd1 net1384 _18292__1384/LO sky130_fd_sc_hd__conb_1
XANTENNA__10216__A1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08290__C1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[20\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13166__A0 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13198__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09007_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[14\]
+ net681 net631 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10615__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09385__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11192__A2 _07092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout686_X net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08312__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12830__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout530 net532 vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09137__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout541 net542 vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__buf_8
Xfanout552 net553 vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__clkbuf_4
X_09909_ _05256_ _05280_ vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__and2_1
Xfanout563 _03692_ vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__buf_1
Xfanout574 net577 vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__buf_2
XANTENNA_fanout853_X net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14330__B net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08345__B1 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12920_ net320 net2831 net474 vssd1 vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__mux2_1
Xfanout596 net597 vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__buf_4
X_12851_ net298 net2779 net481 vssd1 vssd1 vccd1 vccd1 _02783_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_9__f_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_9__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13661__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11802_ _07612_ _07613_ vssd1 vssd1 vccd1 vccd1 _07614_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_4_3__f_wb_clk_i_X clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_68_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15570_ net1281 vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__inv_2
XANTENNA__09845__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12782_ net288 net2453 net489 vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__mux2_1
X_14521_ net1057 vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__inv_2
X_11733_ _07543_ _07544_ vssd1 vssd1 vccd1 vccd1 _07545_ sky130_fd_sc_hd__nor2_1
XFILLER_0_166_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17240_ clknet_leaf_32_wb_clk_i _02870_ _00936_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ net1073 vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__inv_2
X_11664_ net29 net992 _07483_ net1929 vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_25_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13403_ net2640 net232 net419 vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10615_ net2631 net298 net540 vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__mux2_1
X_17171_ clknet_leaf_165_wb_clk_i _02801_ _00867_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14383_ net1528 vssd1 vssd1 vccd1 vccd1 _02993_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11595_ net1606 net1008 net344 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16122_ net1136 vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__inv_2
X_13334_ net244 net2512 net427 vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__mux2_1
X_10546_ _05189_ _05961_ vssd1 vssd1 vccd1 vccd1 _06556_ sky130_fd_sc_hd__xor2_1
XANTENNA__08343__X team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[31\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output183_A net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13157__A0 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16053_ net1173 vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__inv_2
X_18311__1403 vssd1 vssd1 vccd1 vccd1 net1403 _18311__1403/LO sky130_fd_sc_hd__conb_1
X_13265_ net189 net2438 net433 vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_94_Left_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10477_ _06411_ _06490_ net528 vssd1 vssd1 vccd1 vccd1 _06491_ sky130_fd_sc_hd__mux2_1
X_15004_ net1063 vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__inv_2
X_12216_ _08022_ _03510_ vssd1 vssd1 vccd1 vccd1 _03511_ sky130_fd_sc_hd__and2_2
X_13196_ _06216_ net2536 net351 vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__mux2_1
XANTENNA__08584__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08222__C net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12147_ _07950_ _07958_ vssd1 vssd1 vccd1 vccd1 _07959_ sky130_fd_sc_hd__and2_1
XANTENNA__12740__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10930__A2 _06768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12078_ _07874_ _07889_ _07879_ vssd1 vssd1 vccd1 vccd1 _07890_ sky130_fd_sc_hd__a21o_1
X_16955_ clknet_leaf_189_wb_clk_i _02585_ _00651_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11029_ net1045 _07000_ vssd1 vssd1 vccd1 vccd1 _07001_ sky130_fd_sc_hd__nand2_1
X_15906_ net1288 vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__inv_2
X_16886_ clknet_leaf_150_wb_clk_i _02516_ _00582_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15837_ net1269 vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10694__A1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13571__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11880__A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15768_ net1275 vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__inv_2
XANTENNA__09836__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14719_ net1179 vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17507_ clknet_leaf_114_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[10\]
+ _01203_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[10\]
+ sky130_fd_sc_hd__dfrtp_2
X_15699_ net1152 vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__inv_2
X_08240_ net884 net875 net863 vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_99_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17438_ clknet_leaf_67_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[6\]
+ _01134_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08171_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[10\] _04249_
+ vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__nand2_1
X_17369_ clknet_leaf_66_wb_clk_i net1446 _01065_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12915__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_113_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__buf_2
Xoutput122 net122 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__buf_2
XANTENNA__14134__C net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09367__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput133 net133 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__buf_2
Xoutput144 net144 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__clkbuf_4
Xoutput155 net155 vssd1 vssd1 vccd1 vccd1 gpio_out[34] sky130_fd_sc_hd__clkbuf_4
XANTENNA__10906__C1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput166 net166 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__clkbuf_4
XANTENNA__11174__A2 _07101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12371__A1 _03651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08575__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput177 net177 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_56_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput188 net188 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_162_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1019_A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09119__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_68_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__17515__Q team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[18\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08327__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09625_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[2\]
+ net597 _05642_ _05649_ _05650_ vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_69_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13481__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout646_A net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11790__A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09556_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[3\]
+ net682 net644 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05593_ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13623__A1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08507_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[27\]
+ net811 net799 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__a22o_1
X_09487_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[4\]
+ net749 net746 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout434_X net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1176_X net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08438_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[28\]
+ net658 net616 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_156_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08369_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[30\]
+ net830 net769 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout601_X net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12825__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10400_ _06409_ _06417_ _04275_ vssd1 vssd1 vccd1 vccd1 _06418_ sky130_fd_sc_hd__o21a_1
XFILLER_0_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11380_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[0\] _07058_
+ net731 vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10331_ net893 _06347_ _06348_ _06351_ vssd1 vssd1 vccd1 vccd1 _06352_ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10262_ _06003_ _06279_ _06285_ vssd1 vssd1 vccd1 vccd1 _06286_ sky130_fd_sc_hd__o21a_1
XANTENNA__09358__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13050_ net288 net2809 net456 vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11165__A2 _07096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12362__A1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[25\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12001_ net548 _07475_ _07745_ vssd1 vssd1 vccd1 vccd1 _07813_ sky130_fd_sc_hd__nor3_1
XANTENNA__13656__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08566__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12560__S net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10193_ _05913_ _05916_ vssd1 vssd1 vccd1 vccd1 _06219_ sky130_fd_sc_hd__xnor2_4
Xfanout1303 net1311 vssd1 vssd1 vccd1 vccd1 net1303 sky130_fd_sc_hd__clkbuf_4
Xfanout371 net372 vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_108_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16740_ clknet_leaf_183_wb_clk_i _02370_ _00436_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout382 net383 vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__buf_4
X_13952_ _03823_ _03824_ vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__nand2_1
Xfanout393 _03732_ vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12903_ net232 net2458 net474 vssd1 vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__mux2_1
X_16671_ clknet_leaf_153_wb_clk_i _02301_ _00367_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09530__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13883_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[13\]
+ net560 net576 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[13\]
+ net987 vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__a221o_1
XANTENNA__13391__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18410_ net913 vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__clkbuf_1
X_15622_ net1171 vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__inv_2
X_12834_ net242 net2311 net482 vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09818__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18341_ net1330 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
XFILLER_0_29_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18256__Q team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[10\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15553_ net1116 vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12765_ net224 net2602 net490 vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__mux2_1
XANTENNA__09601__C net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14504_ net1223 vssd1 vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18272_ clknet_leaf_36_wb_clk_i _03501_ _01967_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[26\]
+ sky130_fd_sc_hd__dfrtp_4
X_11716_ net356 _07527_ vssd1 vssd1 vccd1 vccd1 _07528_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15484_ net1147 vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12696_ net220 net2615 net498 vssd1 vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17223_ clknet_leaf_199_wb_clk_i _02853_ _00919_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14435_ net1203 vssd1 vssd1 vccd1 vccd1 _00065_ sky130_fd_sc_hd__inv_2
XANTENNA__13917__A2 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12735__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11647_ net16 net989 net916 net1791 vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__o22a_1
XFILLER_0_108_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput13 DAT_I[1] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput24 DAT_I[2] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17154_ clknet_leaf_6_wb_clk_i _02784_ _00850_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09597__A2 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput35 gpio_in[35] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_1
XANTENNA__08254__C1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14366_ _04084_ _04091_ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__nor2_1
Xinput46 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_1
X_11578_ net2927 net1005 _07416_ net357 vssd1 vssd1 vccd1 vccd1 _03335_ sky130_fd_sc_hd__a22o_1
Xinput57 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput68 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__buf_1
X_16105_ net1310 vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold808 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 net2222 sky130_fd_sc_hd__dlygate4sd3_1
X_13317_ net2061 net286 net428 vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__mux2_1
X_10529_ _05829_ _05833_ vssd1 vssd1 vccd1 vccd1 _06540_ sky130_fd_sc_hd__xnor2_4
Xhold819 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2233 sky130_fd_sc_hd__dlygate4sd3_1
X_17085_ clknet_leaf_130_wb_clk_i _02715_ _00781_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_172_Right_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14297_ net381 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_90_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16036_ net1287 vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13248_ net285 net2672 net436 vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13566__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15347__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12470__S _03670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13793__C net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13179_ net285 net2623 net440 vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1508 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net2922 sky130_fd_sc_hd__dlygate4sd3_1
X_17987_ clknet_leaf_64_wb_clk_i _03326_ _01683_ vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18291__1383 vssd1 vssd1 vccd1 vccd1 net1383 _18291__1383/LO sky130_fd_sc_hd__conb_1
Xhold1519 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net2933 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16938_ clknet_leaf_2_wb_clk_i _02568_ _00634_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09521__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16178__A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16869_ clknet_leaf_22_wb_clk_i _02499_ _00565_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_09410_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[6\]
+ net847 net749 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_66_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10938__B _06350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10419__A1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10419__B2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09341_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[7\]
+ net701 net608 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_138_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_186_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_186_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__18393__A net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09272_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[9\]
+ net847 net769 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_62_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_115_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_115_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_74_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08223_ net881 net868 net861 vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14335__A1_N _05256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08154_ net1022 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[5\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[4\] vssd1 vssd1
+ vccd1 vccd1 _04237_ sky130_fd_sc_hd__nand3b_4
XANTENNA__09588__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08796__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08085_ net1026 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__and2b_1
XANTENNA__10165__S _05634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11488__C _07394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1136_A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_951 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12344__A1 _07774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08548__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout596_A net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13476__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12380__S net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1303_A net1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08430__Y _04510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09760__A2 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08987_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[15\]
+ net782 net745 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[15\]
+ _05048_ vssd1 vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout384_X net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout551_X net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout930_A net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout649_X net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08720__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09608_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[2\]
+ net877 net869 net857 vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__and4_1
XFILLER_0_97_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09702__B _05731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10880_ _06791_ _06876_ _06792_ vssd1 vssd1 vccd1 vccd1 _06877_ sky130_fd_sc_hd__a21boi_1
X_18310__1402 vssd1 vssd1 vccd1 vccd1 net1402 _18310__1402/LO sky130_fd_sc_hd__conb_1
XANTENNA__11607__B1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09539_ net570 net533 _05556_ vssd1 vssd1 vccd1 vccd1 _05576_ sky130_fd_sc_hd__o21a_1
XFILLER_0_149_861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout816_X net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_159_Left_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12550_ net1747 _07791_ _03678_ vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11501_ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[11\] _07411_ net1002
+ vssd1 vssd1 vccd1 vccd1 _07412_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12555__S net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12481_ net1683 _07791_ _03673_ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14220_ net728 _04015_ _04016_ vssd1 vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__and3_1
X_11432_ net1050 net1049 vssd1 vssd1 vccd1 vccd1 _07345_ sky130_fd_sc_hd__nor2_4
XFILLER_0_149_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12583__A1 _07789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10043__C1 _06060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14151_ _03800_ net907 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[0\]
+ sky130_fd_sc_hd__nor2_1
X_11363_ _07303_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[1\] net509
+ vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08251__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13102_ net235 net2706 net450 vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10314_ _06282_ _06335_ net520 vssd1 vssd1 vccd1 vccd1 _06336_ sky130_fd_sc_hd__mux2_1
X_14082_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[10\] net980 _03801_
+ vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__o21a_1
XANTENNA__14324__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11294_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[33\] _07097_
+ _07124_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[25\] _07253_
+ vssd1 vssd1 vccd1 vccd1 _07254_ sky130_fd_sc_hd__a221o_1
XANTENNA__08539__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_168_Left_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13386__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17910_ clknet_leaf_76_wb_clk_i _03253_ _01606_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11695__A team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[29\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13033_ net224 net2678 net458 vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__mux2_1
X_10245_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[27\] net906 _06267_
+ _06269_ vssd1 vssd1 vccd1 vccd1 _06270_ sky130_fd_sc_hd__a211o_2
XANTENNA__10346__B1 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11543__C1 team_05_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1100 net1107 vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__clkbuf_2
Xfanout1111 net1127 vssd1 vssd1 vccd1 vccd1 net1111 sky130_fd_sc_hd__buf_4
X_17841_ clknet_leaf_100_wb_clk_i _03184_ _01537_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[87\]
+ sky130_fd_sc_hd__dfrtp_1
X_10176_ net336 _06199_ _06202_ net338 _06194_ vssd1 vssd1 vccd1 vccd1 _06203_ sky130_fd_sc_hd__o221a_1
Xfanout1122 net1127 vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__buf_2
Xfanout1133 net1137 vssd1 vssd1 vccd1 vccd1 net1133 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1144 net1146 vssd1 vssd1 vccd1 vccd1 net1144 sky130_fd_sc_hd__buf_4
Xfanout1155 net1162 vssd1 vssd1 vccd1 vccd1 net1155 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1166 net1175 vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__buf_4
Xfanout1177 net1313 vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__buf_4
X_17772_ clknet_leaf_84_wb_clk_i _03115_ _01468_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_14984_ net1219 vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__inv_2
Xfanout1188 net1190 vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout190 net192 vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__buf_2
Xfanout1199 net1202 vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__buf_4
X_13935_ _03798_ _03809_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[1\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__09503__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16723_ clknet_leaf_165_wb_clk_i _02353_ _00419_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11310__A2 _07113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkload5_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16654_ clknet_leaf_170_wb_clk_i _02284_ _00350_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13866_ net1541 net983 _03769_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[4\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15605_ net1258 vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__inv_2
XFILLER_0_159_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12817_ net288 net2430 net484 vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16585_ clknet_leaf_19_wb_clk_i _02215_ _00281_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13797_ net1578 net975 net725 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[8\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_151_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08228__B net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18324_ net1315 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
X_15536_ net1139 vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__inv_2
X_12748_ net290 net2351 net492 vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18255_ clknet_leaf_41_wb_clk_i _03484_ _01950_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_13_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15467_ net1167 vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__inv_2
XANTENNA__12465__S _03671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12679_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[10\]
+ net339 vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17206_ clknet_leaf_142_wb_clk_i _02836_ _00902_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14418_ net1240 vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18186_ clknet_leaf_42_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[7\]
+ _01881_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15398_ net1280 vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__inv_2
XANTENNA__12574__A1 _07836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08778__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17137_ clknet_leaf_118_wb_clk_i _02767_ _00833_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14349_ _04102_ _04107_ _04121_ vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__or3_1
XANTENNA__08242__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold605 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2019 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold616 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 net2030 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold627 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[9\] vssd1
+ vssd1 vccd1 vccd1 net2041 sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2052 sky130_fd_sc_hd__dlygate4sd3_1
X_17068_ clknet_leaf_0_wb_clk_i _02698_ _00764_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14315__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[19\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold649 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2063 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_51_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13296__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16019_ net1149 vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__inv_2
X_08910_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[16\]
+ net629 net610 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09890_ _04512_ _04554_ _05917_ _04514_ vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__a31o_2
XFILLER_0_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08841_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[18\]
+ net794 net733 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__a22o_1
XANTENNA__18388__A net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1305 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2719 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1316 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 net2730 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1327 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net2741 sky130_fd_sc_hd__dlygate4sd3_1
X_08772_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[19\]
+ net617 net614 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__a22o_1
XANTENNA__10014__A _04818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1338 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2752 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1349 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 net2763 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11301__A2 _07101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08702__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1086_A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09324_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[8\]
+ net820 net792 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[8\]
+ _05371_ vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__a221o_1
XFILLER_0_168_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09255_ net953 _04348_ _04269_ vssd1 vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12375__S _07852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08481__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout609_A _04320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_90_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08206_ _04232_ net962 _04271_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[15\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[16\] vssd1 vssd1
+ vccd1 vccd1 _04289_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_170_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09186_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[10\]
+ net651 net614 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[10\]
+ _05238_ vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_170_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08769__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08137_ _04222_ _04223_ vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__nor2_1
XFILLER_0_133_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10576__B1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_83_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__14306__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[25\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08068_ net1023 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[27\]
+ net970 _04183_ vssd1 vssd1 vccd1 vccd1 _03502_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout880_A net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout599_X net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_12_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12404__A _07840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09194__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10030_ net521 _06058_ vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09733__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout766_X net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08941__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11981_ _07792_ _07787_ _07518_ _07510_ vssd1 vssd1 vccd1 vccd1 _07793_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA_fanout933_X net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11454__S net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13720_ net905 _06408_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[20\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_169_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10932_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[25\] net565 _06922_
+ vssd1 vssd1 vccd1 vccd1 _03431_ sky130_fd_sc_hd__a21o_1
XANTENNA__08329__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13651_ net2443 net319 net390 vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__mux2_1
X_10863_ _06859_ _06818_ _06820_ vssd1 vssd1 vccd1 vccd1 _06860_ sky130_fd_sc_hd__and3b_1
X_12602_ _03605_ net1831 net203 vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__mux2_1
X_16370_ clknet_leaf_125_wb_clk_i _02000_ _00066_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13582_ net2212 net301 net398 vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__mux2_1
X_10794_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[23\] net1040 vssd1
+ vssd1 vccd1 vccd1 _06791_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15321_ net1051 vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__inv_2
X_12533_ net1943 _03605_ net208 vssd1 vssd1 vccd1 vccd1 _03105_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18040_ clknet_leaf_96_wb_clk_i _03378_ _01736_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15252_ net1073 vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__inv_2
X_18290__1382 vssd1 vssd1 vccd1 vccd1 net1382 _18290__1382/LO sky130_fd_sc_hd__conb_1
X_12464_ net1756 _03605_ net212 vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14203_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[7\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[8\]
+ _04003_ vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__and3_1
XANTENNA__11977__X _07789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11415_ _07326_ _07337_ vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__nor2_1
X_15183_ net1281 vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__inv_2
X_12395_ net1671 _03665_ _03660_ vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14134_ team_05_WB.instance_to_wrap.CPU_DAT_O\[17\] net504 net912 vssd1 vssd1 vccd1
+ vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[17\] sky130_fd_sc_hd__and3_1
X_11346_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[11\] net509 net359
+ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[7\] vssd1 vssd1 vccd1
+ vccd1 _03394_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14065_ _03803_ _03868_ _03932_ vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__o21a_1
X_11277_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[106\] _07102_
+ _07115_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[58\] _07214_
+ vssd1 vssd1 vccd1 vccd1 _07238_ sky130_fd_sc_hd__a221o_1
XANTENNA__09185__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13016_ net290 net2886 net460 vssd1 vssd1 vccd1 vccd1 _02625_ sky130_fd_sc_hd__mux2_1
XANTENNA__09724__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10228_ _06016_ _06024_ net526 vssd1 vssd1 vccd1 vccd1 _06253_ sky130_fd_sc_hd__mux2_1
XANTENNA__11531__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_135_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08230__C net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08932__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17824_ clknet_leaf_92_wb_clk_i _03167_ _01520_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instr_fetch vssd1 vssd1
+ vccd1 vccd1 net1416 sky130_fd_sc_hd__dlygate4sd3_1
X_10159_ net893 _06185_ vssd1 vssd1 vccd1 vccd1 _06186_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_85_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17755_ clknet_leaf_77_wb_clk_i _03098_ _01451_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14967_ net1097 vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10769__A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16706_ clknet_leaf_7_wb_clk_i _02336_ _00402_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13918_ net1574 net984 _03795_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[30\]
+ sky130_fd_sc_hd__o21a_1
X_17686_ clknet_leaf_78_wb_clk_i _03029_ _01382_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[124\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14898_ net1239 vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_18_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13849_ net1520 net578 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[27\]
+ sky130_fd_sc_hd__and2_1
X_16637_ clknet_leaf_110_wb_clk_i _02267_ _00333_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_16568_ clknet_leaf_32_wb_clk_i _02198_ _00264_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11598__A2 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08999__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18307_ net1399 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
X_15519_ net1156 vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16499_ clknet_leaf_169_wb_clk_i _02129_ _00195_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09040_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[14\] vssd1
+ vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__inv_2
X_18238_ clknet_leaf_57_wb_clk_i net1514 _01933_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10270__A2 _06293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09948__C1 _05887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18169_ net1038 team_05_WB.instance_to_wrap.total_design.keypad0.next_rows\[1\] _01864_
+ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__dfstp_1
XANTENNA__12923__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08215__A2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold402 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[94\] vssd1 vssd1
+ vccd1 vccd1 net1816 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10009__A _04989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold413 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[43\] vssd1 vssd1
+ vccd1 vccd1 net1827 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_174_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold424 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[55\] vssd1 vssd1
+ vccd1 vccd1 net1838 sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[100\] vssd1 vssd1
+ vccd1 vccd1 net1849 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08261__X _04344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold446 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[54\] vssd1 vssd1
+ vccd1 vccd1 net1860 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold457 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[39\] vssd1 vssd1
+ vccd1 vccd1 net1871 sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 team_05_WB.instance_to_wrap.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1 net1882
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09942_ _05934_ _05969_ _04970_ vssd1 vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__o21bai_1
Xhold479 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[82\] vssd1 vssd1
+ vccd1 vccd1 net1893 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout904 net905 vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__buf_2
XFILLER_0_0_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout915 net183 vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09176__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout926 _04380_ vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__clkbuf_4
X_09873_ _04656_ _04675_ vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__nand2_1
Xfanout937 _04369_ vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__clkbuf_2
Xfanout948 net949 vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_146_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout959 _04244_ vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1102 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2516 sky130_fd_sc_hd__dlygate4sd3_1
X_08824_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[18\]
+ net672 net614 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[18\]
+ _04892_ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__a221o_1
Xhold1113 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2527 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1001_A _07345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1124 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2538 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1135 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net2549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2560 sky130_fd_sc_hd__dlygate4sd3_1
X_08755_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[21\]
+ net847 net775 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__a22o_1
Xhold1157 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2571 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout461_A _03711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1168 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1179 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2593 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08686_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[22\]
+ net700 net646 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_130_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_130_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08149__A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout726_A _03759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout347_X net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11038__A1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_172_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09100__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09307_ _05355_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[8\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_152_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08454__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10261__A2 _06280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09238_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[9\]
+ net635 net616 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[9\]
+ _05286_ vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__a221o_1
XFILLER_0_106_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12538__A1 _03650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09169_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[11\]
+ net771 net741 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[11\]
+ _05222_ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__a221o_1
XANTENNA__12833__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08206__A2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11200_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[46\] _07113_
+ _07116_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[78\] _07151_
+ vssd1 vssd1 vccd1 vccd1 _07165_ sky130_fd_sc_hd__a221o_1
XFILLER_0_161_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12180_ net547 _07690_ vssd1 vssd1 vccd1 vccd1 _07992_ sky130_fd_sc_hd__nand2_4
XANTENNA__12405__Y _03668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14333__B _05801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11131_ _07087_ _07095_ vssd1 vssd1 vccd1 vccd1 _07097_ sky130_fd_sc_hd__nor2_4
XFILLER_0_43_1138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold980 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net2394 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09167__B1 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold991 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net2405 sky130_fd_sc_hd__dlygate4sd3_1
X_11062_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[3\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[4\]
+ _07027_ _07028_ vssd1 vssd1 vccd1 vccd1 _07029_ sky130_fd_sc_hd__and4b_1
XANTENNA__08914__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13664__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10013_ _04778_ net363 _06041_ vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__a21oi_1
X_15870_ net1267 vssd1 vssd1 vccd1 vccd1 _01500_ sky130_fd_sc_hd__inv_2
XANTENNA__10721__B1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input22_A DAT_I[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14821_ net1185 vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_4_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17540_ clknet_leaf_81_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[11\]
+ _01236_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14752_ net1199 vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__inv_2
X_11964_ net501 _07774_ vssd1 vssd1 vccd1 vccd1 _07776_ sky130_fd_sc_hd__or2_1
XANTENNA__08678__C1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13703_ net900 _06706_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[3\]
+ sky130_fd_sc_hd__nor2_1
X_10915_ _06782_ _06783_ vssd1 vssd1 vccd1 vccd1 _06908_ sky130_fd_sc_hd__or2_1
X_17471_ clknet_leaf_40_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[6\]
+ _01167_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_14683_ net1098 vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_80_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08693__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11895_ _07702_ _07703_ _07705_ vssd1 vssd1 vccd1 vccd1 _07707_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_129_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13634_ net1948 net231 net390 vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__mux2_1
X_16422_ clknet_leaf_115_wb_clk_i _02052_ _00118_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10846_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[2\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06843_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16353_ clknet_leaf_149_wb_clk_i _01983_ _00049_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13565_ net2848 net242 net399 vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__mux2_1
X_10777_ _06769_ _06773_ vssd1 vssd1 vccd1 vccd1 _06774_ sky130_fd_sc_hd__nor2_2
XFILLER_0_26_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08445__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15304_ net1223 vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12516_ net1656 _03657_ net209 vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__mux2_1
X_16284_ net1254 vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13496_ net2403 net192 net407 vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__mux2_1
XANTENNA__12529__A1 _03664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18023_ clknet_leaf_96_wb_clk_i _03362_ _01719_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15235_ net1208 vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__inv_2
XANTENNA__08225__C net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12447_ net1742 _03657_ net212 vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__mux2_1
XANTENNA__12743__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14524__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15166_ net1073 vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__inv_2
X_12378_ net1714 _03610_ net216 vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__mux2_1
XANTENNA__10771__B net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14117_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[13\] team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[12\]
+ net978 vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__o21a_1
XANTENNA__10555__A3 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11329_ _04211_ _04215_ vssd1 vssd1 vccd1 vccd1 _07287_ sky130_fd_sc_hd__nor2_1
X_15097_ net1057 vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14048_ _03916_ _03894_ net978 vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13574__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13427__X _03727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15355__A net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17807_ clknet_leaf_90_wb_clk_i _03150_ _01503_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[117\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15999_ net1128 vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08540_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[26\]
+ net817 net789 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[26\]
+ _04615_ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__a221o_1
XFILLER_0_173_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17738_ clknet_leaf_95_wb_clk_i _03081_ _01434_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_141_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08471_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[28\]
+ net843 net780 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[28\]
+ _04549_ vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__a221o_1
X_17669_ clknet_leaf_102_wb_clk_i _03012_ _01365_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[107\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12918__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08436__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_114_Left_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11440__A1 _07349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09023_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[14\]
+ net817 net740 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout307_A net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1049_A team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold210 team_05_WB.instance_to_wrap.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 net1624
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold221 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[69\] vssd1 vssd1
+ vccd1 vccd1 net1635 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold232 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[20\] vssd1 vssd1
+ vccd1 vccd1 net1646 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17518__Q team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[21\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold243 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[36\] vssd1 vssd1
+ vccd1 vccd1 net1657 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[45\] vssd1 vssd1
+ vccd1 vccd1 net1668 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold265 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[120\] vssd1 vssd1
+ vccd1 vccd1 net1679 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10026__X _06055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold276 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[98\] vssd1 vssd1
+ vccd1 vccd1 net1690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[18\] vssd1 vssd1
+ vccd1 vccd1 net1701 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09149__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout701 _04293_ vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__buf_4
Xhold298 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[56\] vssd1 vssd1
+ vccd1 vccd1 net1712 sky130_fd_sc_hd__dlygate4sd3_1
X_09925_ _05812_ _05952_ _05810_ vssd1 vssd1 vccd1 vccd1 _05954_ sky130_fd_sc_hd__a21o_1
Xfanout712 _04288_ vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__buf_2
XFILLER_0_102_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout723 net724 vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_165_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout734 net736 vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_123_Left_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout676_A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13484__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout745 _04417_ vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__buf_6
XANTENNA__15265__A net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout756 net759 vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__buf_6
X_09856_ _04818_ _04838_ vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__or2_1
Xfanout767 _04408_ vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__buf_4
Xfanout778 net781 vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10703__B1 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout789 _04400_ vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__buf_4
X_08807_ net853 _04865_ _04866_ _04876_ vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__or4_1
XFILLER_0_147_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09787_ net349 _05329_ vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__nand2_1
Xclkbuf_4_8__f_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_8__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_fanout464_X net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout843_A net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08738_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[21\]
+ net701 net669 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[21\]
+ _04809_ vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__a221o_1
XFILLER_0_68_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09321__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08669_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[23\]
+ net766 net749 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[23\]
+ _04742_ vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout631_X net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08675__A2 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10700_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[3\] team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[2\]
+ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[4\] vssd1 vssd1 vccd1
+ vccd1 _06702_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09710__B net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11680_ net66 net65 net68 net67 vssd1 vssd1 vccd1 vccd1 _07494_ sky130_fd_sc_hd__or4_1
XFILLER_0_95_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14328__B _05596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10631_ _04174_ net902 net897 _06636_ _06634_ vssd1 vssd1 vccd1 vccd1 _06637_ sky130_fd_sc_hd__o221a_4
XANTENNA__08427__A2 _04366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08326__B net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13350_ net286 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[10\]
+ net425 vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10562_ net2083 net279 net539 vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12301_ _03594_ _03595_ _03512_ vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13659__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12563__S _03678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13281_ net282 net2139 net433 vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10493_ _06430_ _06505_ net532 vssd1 vssd1 vccd1 vccd1 _06506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09388__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15020_ net1109 vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__inv_2
X_12232_ _08014_ _08018_ _03525_ vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_20_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14063__B net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12163_ _07920_ _07962_ _07969_ vssd1 vssd1 vccd1 vccd1 _07975_ sky130_fd_sc_hd__and3_1
XFILLER_0_102_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11114_ _07078_ _07079_ vssd1 vssd1 vccd1 vccd1 _07081_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_9_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16971_ clknet_leaf_186_wb_clk_i _02601_ _00667_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_12094_ _07895_ _07897_ _07900_ vssd1 vssd1 vccd1 vccd1 _07906_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15922_ net1296 vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__inv_2
X_11045_ _07014_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[4\] net569
+ vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__mux2_1
XANTENNA__09444__Y team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[5\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18259__Q team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15853_ net1257 vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__inv_2
XANTENNA__09604__C net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14804_ net1066 vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__inv_2
X_15784_ net1257 vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__inv_2
X_12996_ net199 net2559 net462 vssd1 vssd1 vccd1 vccd1 _02645_ sky130_fd_sc_hd__mux2_1
XANTENNA__09312__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09901__A net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17523_ clknet_leaf_73_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[26\]
+ _01219_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[26\]
+ sky130_fd_sc_hd__dfrtp_2
X_11947_ _07734_ _07736_ _07730_ vssd1 vssd1 vccd1 vccd1 _07759_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14735_ net1239 vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__inv_2
XANTENNA__12738__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08666__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17454_ clknet_leaf_57_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[22\]
+ _01150_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_14666_ net1121 vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__inv_2
XANTENNA__10473__A2 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11878_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[3\] net993 vssd1
+ vssd1 vccd1 vccd1 _07690_ sky130_fd_sc_hd__nand2_2
XANTENNA__08517__A _04573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13617_ net2197 net302 net394 vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__mux2_1
X_16405_ clknet_leaf_175_wb_clk_i _02035_ _00101_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10829_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[9\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06826_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17385_ clknet_leaf_49_wb_clk_i net1417 _01081_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14597_ net1191 vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__inv_2
XANTENNA__08418__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08236__B net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16336_ net1117 vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__inv_2
X_13548_ net2279 net288 net400 vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__mux2_1
XANTENNA__09091__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13569__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11878__A team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16267_ net1123 vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_97_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13479_ net283 net2638 net409 vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13796__C net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14372__A0 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18006_ clknet_leaf_62_wb_clk_i _03345_ _01702_ vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09379__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15218_ net1235 vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16198_ net1146 vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11186__B1 _07121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1036 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_93_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15149_ net1080 vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09710_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[0\]
+ net944 net936 net926 vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_143_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09354__Y team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09551__B1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09641_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[1\]
+ net940 net935 net932 vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_160_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09572_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[2\]
+ net940 net932 net930 vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__and4_1
XANTENNA__08106__A1 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08523_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[26\]
+ net709 net627 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[26\]
+ _04599_ vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_69_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08657__A2 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout257_A _06442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10464__A2 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08454_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[28\]
+ net718 _04529_ _04532_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__o22a_2
XFILLER_0_77_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08385_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[30\]
+ net592 _04456_ _04465_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[30\]
+ sky130_fd_sc_hd__o22a_4
XFILLER_0_135_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout424_A _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1166_A net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12610__A0 _03623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09082__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13479__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11788__A team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout212_X net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12383__S net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11140__X _07106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09006_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[14\]
+ net669 net654 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[14\]
+ _05066_ vssd1 vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_167_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11177__B1 _07124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10924__A0 _06273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_131_Left_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout960_A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout581_X net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout520 net522 vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout679_X net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout531 net532 vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__buf_2
Xfanout542 _04260_ vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__buf_4
X_09908_ _05165_ _05185_ vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__and2b_1
Xfanout553 _06052_ vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09705__B net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout564 net567 vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__clkbuf_4
Xfanout575 net576 vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__buf_2
XANTENNA__09542__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09839_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[20\]
+ net760 net756 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__a22o_1
Xfanout597 _04323_ vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout846_X net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08896__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12429__A0 _03605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12850_ net287 net2509 net480 vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__mux2_1
X_11801_ _07589_ _07596_ _07593_ vssd1 vssd1 vccd1 vccd1 _07613_ sky130_fd_sc_hd__a21o_1
XANTENNA__12558__S net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12781_ net292 net2577 net488 vssd1 vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__mux2_1
Xclkbuf_3_1_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08648__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11462__S net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_140_Left_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14520_ net1242 vssd1 vssd1 vccd1 vccd1 _00150_ sky130_fd_sc_hd__inv_2
X_11732_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[11\] net550 net998
+ _07525_ vssd1 vssd1 vccd1 vccd1 _07544_ sky130_fd_sc_hd__and4_1
XANTENNA__08337__A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14451_ net1212 vssd1 vssd1 vccd1 vccd1 _00081_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11663_ net30 net990 net917 net1882 vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__o22a_1
XFILLER_0_166_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_153_Right_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ net1951 net235 net418 vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__mux2_1
X_10614_ _06618_ _06620_ _04264_ vssd1 vssd1 vccd1 vccd1 _06621_ sky130_fd_sc_hd__a21oi_4
XANTENNA__10207__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17170_ clknet_leaf_127_wb_clk_i _02800_ _00866_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_14382_ net1517 vssd1 vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11594_ net131 net1011 net346 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09073__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16121_ net1136 vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__inv_2
XANTENNA__13389__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11698__A team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[24\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13333_ net222 net2195 net426 vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08281__B1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[24\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10545_ net1941 net284 net542 vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08820__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16052_ net1173 vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13264_ net193 net2467 net435 vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10476_ _06447_ _06489_ net518 vssd1 vssd1 vccd1 vccd1 _06490_ sky130_fd_sc_hd__mux2_1
XANTENNA__11168__B1 _07126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15003_ net1098 vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__inv_2
XANTENNA__11985__X _07797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12215_ _07867_ _07894_ _03509_ _07552_ vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__or4b_4
XFILLER_0_122_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13195_ net193 net2528 net352 vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12146_ _07902_ _07910_ _07952_ _07955_ _07956_ vssd1 vssd1 vccd1 vccd1 _07958_ sky130_fd_sc_hd__a32o_1
XANTENNA__10391__A1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12077_ _07865_ _07876_ _07869_ vssd1 vssd1 vccd1 vccd1 _07889_ sky130_fd_sc_hd__a21o_1
X_16954_ clknet_leaf_31_wb_clk_i _02584_ _00650_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09533__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15905_ net1295 vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__inv_2
X_11028_ _06830_ _06831_ _06850_ vssd1 vssd1 vccd1 vccd1 _07000_ sky130_fd_sc_hd__a21o_1
X_16885_ clknet_leaf_71_wb_clk_i _02515_ _00581_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08887__A2 _04383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15836_ net1293 vssd1 vssd1 vccd1 vccd1 _01466_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13093__A0 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11880__B _07690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12468__S _03670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10777__A _06769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15767_ net1302 vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__inv_2
X_12979_ net272 net2663 net464 vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__mux2_1
XANTENNA__08639__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17506_ clknet_leaf_110_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[9\]
+ _01202_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_14718_ net1062 vssd1 vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15698_ net1152 vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__inv_2
XANTENNA__10496__B net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17437_ clknet_leaf_67_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[5\]
+ _01133_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_14649_ net1057 vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08170_ _04252_ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__inv_2
X_17368_ clknet_leaf_60_wb_clk_i net1440 _01064_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09064__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10603__C1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13299__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16319_ net1141 vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17299_ clknet_leaf_166_wb_clk_i _02929_ _00995_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput123 net123 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_140_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12931__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput134 net134 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__buf_2
Xoutput145 net145 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__clkbuf_4
XANTENNA__14712__A net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput156 net156 vssd1 vssd1 vccd1 vccd1 gpio_out[35] sky130_fd_sc_hd__clkbuf_4
XANTENNA__10906__B1 _06898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput167 net167 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_110_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput178 net178 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_162_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13328__A team_05_WB.instance_to_wrap.total_design.core.instr_fetch vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09524__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10134__A1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09624_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[2\]
+ net707 _05636_ _05644_ _05647_ vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_108_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09555_ _05586_ _05588_ _05589_ _05591_ vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__or4_1
XANTENNA__12378__S net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_37_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout541_A net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout639_A _04312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1283_A net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11135__X _07101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08506_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[27\]
+ net819 net807 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[27\]
+ _04583_ vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__a221o_1
XFILLER_0_144_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09486_ _05519_ _05521_ _05523_ _05525_ vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__or4_1
XFILLER_0_109_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08437_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[28\]
+ net696 net641 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[28\]
+ _04515_ vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__a221o_1
XFILLER_0_110_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout806_A net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout427_X net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08368_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[30\]
+ net842 net811 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[30\]
+ _04448_ vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__a221o_1
XFILLER_0_34_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09055__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08263__B1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[31\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08802__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08299_ net948 net1014 net926 vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__and3_1
XANTENNA__09460__C1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13002__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10330_ net890 _06350_ vssd1 vssd1 vccd1 vccd1 _06351_ sky130_fd_sc_hd__and2_1
XFILLER_0_131_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout796_X net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10261_ net338 _06280_ _06284_ net336 _06281_ vssd1 vssd1 vccd1 vccd1 _06285_ sky130_fd_sc_hd__o221a_1
XANTENNA__12841__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12000_ _07477_ _07517_ _07796_ vssd1 vssd1 vccd1 vccd1 _07812_ sky130_fd_sc_hd__a21oi_4
X_10192_ _05916_ _05994_ vssd1 vssd1 vccd1 vccd1 _06218_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout963_X net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1304 net1306 vssd1 vssd1 vccd1 vccd1 net1304 sky130_fd_sc_hd__buf_4
Xfanout350 _03717_ vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__buf_6
Xfanout361 net362 vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__buf_2
Xfanout372 _05576_ vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__clkbuf_4
X_13951_ _03821_ _03822_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__a21o_1
Xfanout383 _04265_ vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__buf_6
XANTENNA__11322__B1 _07110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout394 net395 vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__buf_6
XANTENNA__08869__A2 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13672__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12902_ net235 net2394 net474 vssd1 vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__mux2_1
X_13882_ net1557 net982 _03777_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[12\]
+ sky130_fd_sc_hd__o21a_1
X_16670_ clknet_leaf_184_wb_clk_i _02300_ _00366_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_15621_ net1169 vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__inv_2
X_12833_ net223 net2489 net481 vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_1062 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18340_ net1329 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
XFILLER_0_5_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15552_ net1117 vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__inv_2
X_12764_ net221 net2917 net491 vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09294__A2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09601__D net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11715_ _07519_ _07521_ _07526_ vssd1 vssd1 vccd1 vccd1 _07527_ sky130_fd_sc_hd__or3b_2
XFILLER_0_56_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14503_ net1104 vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__inv_2
X_15483_ net1147 vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__inv_2
X_18271_ clknet_leaf_36_wb_clk_i _03500_ _01966_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[25\]
+ sky130_fd_sc_hd__dfrtp_4
X_12695_ net190 net2745 net498 vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13701__A net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17222_ clknet_leaf_119_wb_clk_i _02852_ _00918_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14434_ net1217 vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_42_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11646_ net17 net989 net916 net2797 vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__o22a_1
XANTENNA__09046__A2 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18272__Q team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[26\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput14 DAT_I[20] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17153_ clknet_leaf_148_wb_clk_i _02783_ _00849_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_14365_ _04087_ _04137_ _04092_ vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__o21ba_1
Xinput25 DAT_I[30] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
Xinput36 gpio_in[36] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_1
X_11577_ net2086 net1005 _07412_ net357 vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__a22o_1
Xinput47 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput58 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__buf_1
X_16104_ net1300 vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13316_ net2046 net292 net428 vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14327__B1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput69 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_1
X_10528_ _05833_ _05962_ _06538_ vssd1 vssd1 vccd1 vccd1 _06539_ sky130_fd_sc_hd__a21oi_1
X_17084_ clknet_leaf_165_wb_clk_i _02714_ _00780_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold809 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2223 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14296_ _04065_ _04067_ _04068_ vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__and3_1
XFILLER_0_161_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08233__C net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_41_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16035_ net1287 vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13247_ net274 net2242 net438 vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_90_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10459_ net337 _06299_ _06470_ net348 _06473_ vssd1 vssd1 vccd1 vccd1 _06474_ sky130_fd_sc_hd__o221a_1
XFILLER_0_62_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12751__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13178_ net275 net2794 net442 vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__mux2_1
XANTENNA__10364__A1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12129_ _07936_ _07940_ _07931_ vssd1 vssd1 vccd1 vccd1 _07941_ sky130_fd_sc_hd__a21o_1
XANTENNA__10271__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17986_ clknet_leaf_63_wb_clk_i _03325_ _01682_ vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__dfrtp_2
Xhold1509 net164 vssd1 vssd1 vccd1 vccd1 net2923 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09506__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16937_ clknet_leaf_14_wb_clk_i _02567_ _00633_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11313__B1 _07111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13582__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16868_ clknet_leaf_182_wb_clk_i _02498_ _00564_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15819_ net1305 vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__inv_2
X_16799_ clknet_leaf_153_wb_clk_i _02429_ _00495_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09340_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[7\]
+ net692 net684 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[7\]
+ _05386_ vssd1 vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09285__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09271_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[9\]
+ net819 net807 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[9\]
+ _05320_ vssd1 vssd1 vccd1 vccd1 _05321_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_103_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08493__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12926__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14707__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08222_ net878 net867 net863 vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__and3_4
XANTENNA_clkbuf_leaf_80_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08705__A _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09037__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08153_ net1022 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[5\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[4\] vssd1 vssd1
+ vccd1 vccd1 _04236_ sky130_fd_sc_hd__and3b_2
XANTENNA__12041__A1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[19\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08245__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_155_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_155_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_16_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_151_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14145__C net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14318__B1 _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10052__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08084_ net1024 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[19\]
+ net973 _04191_ vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1031_A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13541__A1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10355__A1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10355__B2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout491_A _03700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17526__Q team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[29\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08986_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[15\]
+ net798 net760 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout756_A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13492__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_127_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09607_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[2\]
+ net886 net868 _04296_ vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_27_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout923_A _05213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11607__A1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[18\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09538_ net533 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[3\]
+ sky130_fd_sc_hd__inv_2
XANTENNA__11607__B2 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10210__A _05634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09276__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09469_ _04246_ net1017 _04233_ net958 vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__o211a_1
XANTENNA__08484__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout711_X net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12836__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout809_X net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11500_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[11\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[11\]
+ net1034 vssd1 vssd1 vccd1 vccd1 _07411_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12480_ net1899 _07789_ _03673_ vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09028__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11431_ team_05_WB.instance_to_wrap.wishbone.curr_state\[2\] team_05_WB.instance_to_wrap.wishbone.curr_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _07344_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14150_ _03685_ team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.next_next_data_read
+ team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.next_next_fetch vssd1 vssd1
+ vccd1 vccd1 _03994_ sky130_fd_sc_hd__or3b_2
X_11362_ _07289_ _07298_ _07302_ _07291_ _07301_ vssd1 vssd1 vccd1 vccd1 _07303_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13101_ net238 net2089 net451 vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13667__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10313_ _06165_ _06167_ vssd1 vssd1 vccd1 vccd1 _06335_ sky130_fd_sc_hd__nand2_1
XANTENNA__12571__S _03678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14081_ net910 _03948_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[8\]
+ sky130_fd_sc_hd__nor2_1
X_11293_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[105\] _07102_
+ _07103_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[113\] _07252_
+ vssd1 vssd1 vccd1 vccd1 _07253_ sky130_fd_sc_hd__a221o_1
XFILLER_0_131_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13032_ net219 net2321 net458 vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__mux2_1
XANTENNA_input52_A wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10244_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[27\] net968
+ _04247_ _06268_ vssd1 vssd1 vccd1 vccd1 _06269_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09200__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11543__B1 _07349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1101 net1103 vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__buf_4
X_17840_ clknet_leaf_104_wb_clk_i _03183_ _01536_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[86\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1112 net1120 vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__buf_4
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_125_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10175_ _06200_ _06201_ net528 vssd1 vssd1 vccd1 vccd1 _06202_ sky130_fd_sc_hd__mux2_1
Xfanout1123 net1126 vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__buf_4
Xfanout1134 net1137 vssd1 vssd1 vccd1 vccd1 net1134 sky130_fd_sc_hd__buf_4
Xfanout1145 net1146 vssd1 vssd1 vccd1 vccd1 net1145 sky130_fd_sc_hd__buf_4
Xfanout1156 net1162 vssd1 vssd1 vccd1 vccd1 net1156 sky130_fd_sc_hd__buf_4
Xfanout1167 net1170 vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__buf_4
XFILLER_0_156_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17771_ clknet_leaf_90_wb_clk_i _03114_ _01467_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14983_ net1105 vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__inv_2
Xfanout1178 net1181 vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__buf_4
Xfanout1189 net1190 vssd1 vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__buf_4
Xfanout191 net192 vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__clkbuf_2
X_16722_ clknet_leaf_123_wb_clk_i _02352_ _00418_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13934_ team_05_WB.instance_to_wrap.CPU_DAT_O\[1\] net506 _03808_ vssd1 vssd1 vccd1
+ vccd1 _03809_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_1112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09181__A net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18267__Q team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[21\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16653_ clknet_leaf_161_wb_clk_i _02283_ _00349_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13865_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[4\]
+ net559 net575 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[4\]
+ net986 vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09612__C net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_69_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15604_ net1259 vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__inv_2
X_12816_ net291 net2677 net484 vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16584_ clknet_leaf_204_wb_clk_i _02214_ _00280_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13796_ net1602 net976 net725 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[7\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__09267__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18323_ net1314 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_29_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08228__C net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15535_ net1140 vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__inv_2
X_12747_ net278 net2397 net492 vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__mux2_1
XANTENNA__12746__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11503__X _07414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18254_ clknet_leaf_40_wb_clk_i _03483_ _01949_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_15466_ net1158 vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__inv_2
X_12678_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[11\]
+ net339 vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_13_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17205_ clknet_leaf_23_wb_clk_i _02835_ _00901_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_14417_ net1212 vssd1 vssd1 vccd1 vccd1 _00047_ sky130_fd_sc_hd__inv_2
X_11629_ net2697 net1008 net345 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__a22o_1
X_18185_ clknet_leaf_40_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[6\]
+ _01880_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15397_ net1196 vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17136_ clknet_leaf_137_wb_clk_i _02766_ _00832_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_164_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14348_ _05078_ _05099_ _04093_ _04115_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__a211o_1
XANTENNA__10585__A1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold606 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2020 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold617 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2031 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13577__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15358__A net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold628 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net2042 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold639 net101 vssd1 vssd1 vccd1 vccd1 net2053 sky130_fd_sc_hd__dlygate4sd3_1
X_14279_ _06706_ _06729_ _06743_ _06756_ vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__and4_1
XANTENNA__12481__S _03673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17067_ clknet_leaf_188_wb_clk_i _02697_ _00763_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_59_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16018_ net1143 vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08840_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[18\]
+ net756 net745 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[18\]
+ _04906_ vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_55_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1034 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1306 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2720 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1317 team_05_WB.instance_to_wrap.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 net2731
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08771_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[19\]
+ net683 net624 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__a22o_1
Xhold1328 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net2742 sky130_fd_sc_hd__dlygate4sd3_1
X_17969_ clknet_leaf_106_wb_clk_i _03308_ _01665_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__dfrtp_1
Xhold1339 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2753 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09323_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[8\]
+ _04366_ net766 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[8\]
+ net856 vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__a221o_1
XFILLER_0_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08466__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12509__X _03676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09254_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[9\]
+ net717 _05304_ vssd1 vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__o21ai_4
XANTENNA_fanout1079_A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08435__A _04490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08205_ net884 net874 net870 vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__and3_4
XFILLER_0_141_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12014__A1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[31\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13211__A0 _06536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09185_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[10\]
+ net659 net617 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08136_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[3\] team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[2\]
+ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[1\] team_05_WB.instance_to_wrap.total_design.data_from_keypad\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__or4b_1
XFILLER_0_133_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09430__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13487__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12391__S _07852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08067_ net1023 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__and2b_1
XANTENNA__09537__Y _05575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1034_X net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_15__f_wb_clk_i_X clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout494_X net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_52_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout661_X net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08969_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[15\]
+ net664 net644 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[15\]
+ _05031_ vssd1 vssd1 vccd1 vccd1 _05032_ sky130_fd_sc_hd__a221o_1
XANTENNA__17633__D team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout759_X net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11980_ net501 _07714_ vssd1 vssd1 vccd1 vccd1 _07792_ sky130_fd_sc_hd__nor2_1
XANTENNA__09713__B net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09497__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10931_ net960 _06918_ _06921_ vssd1 vssd1 vccd1 vccd1 _06922_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10211__Y _06237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10500__A1 _06033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout926_X net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18369__1354 vssd1 vssd1 vccd1 vccd1 _18369__1354/HI net1354 sky130_fd_sc_hd__conb_1
XANTENNA__10500__B2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08329__B net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10862_ _06824_ _06825_ _06855_ _06822_ _06821_ vssd1 vssd1 vccd1 vccd1 _06859_ sky130_fd_sc_hd__o311a_1
X_13650_ net2800 net302 net390 vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12601_ net1659 _07797_ _03680_ vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13581_ net2257 net288 net397 vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__mux2_1
XANTENNA__08457__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12566__S _03678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10793_ _06788_ _06789_ vssd1 vssd1 vccd1 vccd1 _06790_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12532_ _07797_ net1770 _03675_ vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__mux2_1
XANTENNA__10264__B1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15320_ net1244 vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12463_ net1641 _07797_ _03670_ vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__mux2_1
X_15251_ net1214 vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14202_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[7\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[6\]
+ _04000_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[8\] vssd1
+ vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__a31o_1
X_11414_ net2041 _07325_ vssd1 vssd1 vccd1 vccd1 _07337_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15182_ net1180 vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__inv_2
X_12394_ _07864_ net355 vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__and2_2
XFILLER_0_34_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14133_ net2971 net502 net911 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[16\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__13397__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11345_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[12\] net509 net359
+ net980 vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14064_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[15\] net978 team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[13\]
+ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[12\] vssd1 vssd1 vccd1
+ vccd1 _03932_ sky130_fd_sc_hd__or4_1
XFILLER_0_123_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11276_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[50\] _07117_
+ _07118_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[66\] _07236_
+ vssd1 vssd1 vccd1 vccd1 _07237_ sky130_fd_sc_hd__a221o_1
XANTENNA__10319__A1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_59 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09607__C net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_18_Left_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13015_ net278 net2427 net460 vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__mux2_1
X_10227_ net525 _06009_ vssd1 vssd1 vccd1 vccd1 _06252_ sky130_fd_sc_hd__or2_1
XANTENNA__14810__A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10115__A _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09463__X team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[5\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17823_ clknet_leaf_87_wb_clk_i _03166_ _01519_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09904__A _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08932__B2 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10158_ _05918_ _05927_ vssd1 vssd1 vccd1 vccd1 _06185_ sky130_fd_sc_hd__xnor2_4
XTAP_TAPCELL_ROW_33_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[17\]
+ vssd1 vssd1 vccd1 vccd1 net1417 sky130_fd_sc_hd__dlygate4sd3_1
X_17754_ clknet_leaf_102_wb_clk_i _03097_ _01450_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14966_ net1084 vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_85_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10089_ _06116_ vssd1 vssd1 vccd1 vccd1 _06117_ sky130_fd_sc_hd__inv_2
XANTENNA__09488__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10769__B _06766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16705_ clknet_leaf_149_wb_clk_i _02335_ _00401_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13917_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[30\]
+ net561 net574 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[30\]
+ net985 vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__a221o_1
XFILLER_0_159_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11295__A2 _07119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17685_ clknet_leaf_103_wb_clk_i _03028_ _01381_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[123\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12492__A1 _03645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08696__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14897_ net1192 vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08239__B net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16636_ clknet_leaf_155_wb_clk_i _02266_ _00332_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13848_ net1530 net579 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[26\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08448__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12476__S net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16567_ clknet_leaf_143_wb_clk_i _02197_ _00263_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13779_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[29\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[28\] team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[31\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[30\] vssd1
+ vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__or4_1
XANTENNA__13799__C net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11380__S net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18306_ net1398 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
XFILLER_0_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15518_ net1148 vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16498_ clknet_leaf_126_wb_clk_i _02128_ _00194_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09660__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18237_ clknet_leaf_57_wb_clk_i net1479 _01932_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15449_ net1168 vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18168_ net1038 team_05_WB.instance_to_wrap.total_design.keypad0.next_rows\[0\] _01863_
+ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09412__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold403 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[44\] vssd1 vssd1
+ vccd1 vccd1 net1817 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_3_3_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold414 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[121\] vssd1 vssd1
+ vccd1 vccd1 net1828 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17119_ clknet_leaf_156_wb_clk_i _02749_ _00815_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold425 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[113\] vssd1 vssd1
+ vccd1 vccd1 net1839 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08620__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold436 net94 vssd1 vssd1 vccd1 vccd1 net1850 sky130_fd_sc_hd__dlygate4sd3_1
X_18099_ clknet_leaf_53_wb_clk_i _03422_ _01795_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_40_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold447 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[81\] vssd1 vssd1
+ vccd1 vccd1 net1861 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13100__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold458 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[60\] vssd1 vssd1
+ vccd1 vccd1 net1872 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold469 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[1\] vssd1 vssd1
+ vccd1 vccd1 net1883 sky130_fd_sc_hd__dlygate4sd3_1
X_09941_ _05934_ _05969_ vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_129_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18399__A net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout905 net906 vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__clkbuf_4
Xfanout916 _07484_ vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__buf_2
XFILLER_0_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout927 net929 vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__buf_2
X_09872_ _04656_ _04675_ vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__nor2_1
XANTENNA__10025__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout938 net939 vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__buf_2
Xfanout949 _04363_ vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_146_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09373__X team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1103 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2517 sky130_fd_sc_hd__dlygate4sd3_1
X_08823_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[18\]
+ net660 net636 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_146_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1114 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2528 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10730__A1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_7__f_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_7__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_31_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout287_A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1125 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net2539 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1136 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net2550 sky130_fd_sc_hd__dlygate4sd3_1
X_08754_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[21\]
+ net834 net742 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[21\]
+ _04825_ vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__a221o_1
Xhold1147 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net2561 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1158 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 net2572 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09479__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1169 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net2583 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11286__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12483__A1 _07793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08685_ _04757_ vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__inv_2
XANTENNA__08687__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10031__Y _06060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout454_A _03713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08439__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_170_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_170_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_48_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout621_A net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09306_ _04246_ _04351_ _05352_ _05353_ vssd1 vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout719_A _04285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08165__A net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09237_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[9\]
+ net680 net645 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[9\]
+ _05287_ vssd1 vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1151_X net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout507_X net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09168_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[11\]
+ net829 net768 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_118_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09403__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08119_ net1028 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__and2b_1
XANTENNA__11210__A2 _07102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09099_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[12\]
+ net687 net601 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08611__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09708__B net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13010__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11130_ _07039_ _07095_ vssd1 vssd1 vccd1 vccd1 _07096_ sky130_fd_sc_hd__nor2_4
Xhold970 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2395 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout876_X net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11061_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[5\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[14\]
+ vssd1 vssd1 vccd1 vccd1 _07028_ sky130_fd_sc_hd__nor2_1
Xhold992 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net2406 sky130_fd_sc_hd__dlygate4sd3_1
X_10012_ net378 net363 vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__nor2_1
XANTENNA__10721__A1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11465__S net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14820_ net1205 vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__inv_2
XANTENNA__11692__C net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input15_A DAT_I[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11277__A2 _07102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14751_ net1184 vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11963_ net501 _07774_ vssd1 vssd1 vccd1 vccd1 _07775_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13680__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13702_ net900 _06729_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[2\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__10485__B1 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17470_ clknet_leaf_38_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[5\]
+ _01166_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10914_ _05912_ _06906_ vssd1 vssd1 vccd1 vccd1 _06907_ sky130_fd_sc_hd__nand2_2
X_14682_ net1055 vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11894_ _07705_ vssd1 vssd1 vccd1 vccd1 _07706_ sky130_fd_sc_hd__inv_2
XFILLER_0_168_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16421_ clknet_leaf_180_wb_clk_i _02051_ _00117_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10845_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[0\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[0\]
+ _06840_ _06838_ vssd1 vssd1 vccd1 vccd1 _06842_ sky130_fd_sc_hd__a31o_1
X_13633_ net2579 net234 net390 vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16352_ clknet_leaf_132_wb_clk_i _01982_ _00048_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10776_ team_05_WB.instance_to_wrap.total_design.core.data_access team_05_WB.instance_to_wrap.total_design.core.disable_pc_reg
+ _06772_ team_05_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 _06773_ sky130_fd_sc_hd__and4bb_1
X_13564_ net2010 net223 net398 vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15303_ net1106 vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__inv_2
X_12515_ _07791_ net1824 _03675_ vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__mux2_1
X_16283_ net1254 vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__inv_2
X_13495_ net2179 net194 net405 vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__mux2_1
XANTENNA__08850__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18022_ clknet_leaf_96_wb_clk_i _03361_ _01718_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12446_ net1767 _07791_ _03670_ vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__mux2_1
X_15234_ net1193 vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__inv_2
XANTENNA__11201__A2 _07123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12377_ net1652 _03655_ net217 vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15165_ net1088 vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_26_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11328_ net34 net35 net37 net36 vssd1 vssd1 vccd1 vccd1 _07286_ sky130_fd_sc_hd__or4b_2
X_14116_ net910 _03980_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[11\]
+ sky130_fd_sc_hd__nor2_1
X_15096_ net1201 vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15636__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14047_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[12\] _03893_ _03894_
+ vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__a21bo_1
X_11259_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[99\] _07123_
+ _07126_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[83\] _07220_
+ vssd1 vssd1 vccd1 vccd1 _07221_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12612__X _03683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14540__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17806_ clknet_leaf_81_wb_clk_i _03149_ _01502_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[116\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08381__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15998_ net1130 vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_167_Right_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17737_ clknet_leaf_100_wb_clk_i _03080_ _01433_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11268__A2 _07125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14949_ net1191 vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__inv_2
XANTENNA__08669__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Left_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13590__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08470_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[28\]
+ net792 net743 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17668_ clknet_leaf_93_wb_clk_i _03011_ _01364_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16619_ clknet_leaf_185_wb_clk_i _02249_ _00315_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17599_ clknet_leaf_80_wb_clk_i _02970_ _01295_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09094__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11440__A2 _07351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12934__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08841__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09022_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[14\]
+ net851 net773 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[14\]
+ _05081_ vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold200 team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.state\[0\] vssd1 vssd1
+ vccd1 vccd1 net1614 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold211 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[106\] vssd1 vssd1
+ vccd1 vccd1 net1625 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout202_A _03683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold222 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[79\] vssd1 vssd1
+ vccd1 vccd1 net1636 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold233 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[3\] vssd1 vssd1
+ vccd1 vccd1 net1647 sky130_fd_sc_hd__dlygate4sd3_1
X_18368__1353 vssd1 vssd1 vccd1 vccd1 _18368__1353/HI net1353 sky130_fd_sc_hd__conb_1
Xhold244 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[74\] vssd1 vssd1
+ vccd1 vccd1 net1658 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10400__B1 _04275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold255 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[105\] vssd1 vssd1
+ vccd1 vccd1 net1669 sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[59\] vssd1 vssd1
+ vccd1 vccd1 net1680 sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[110\] vssd1 vssd1
+ vccd1 vccd1 net1691 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold288 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[37\] vssd1 vssd1
+ vccd1 vccd1 net1702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[92\] vssd1 vssd1
+ vccd1 vccd1 net1713 sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ _05812_ _05952_ vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout702 _04293_ vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__buf_2
Xfanout713 _04288_ vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_165_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout724 net726 vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__buf_2
XFILLER_0_0_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1111_A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout735 net736 vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_165_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout746 net747 vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__clkbuf_8
X_09855_ _05883_ vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__inv_2
Xfanout757 net759 vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__clkbuf_8
XANTENNA_input7_A DAT_I[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout571_A net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout768 net770 vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__buf_6
Xfanout779 net781 vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08372__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout669_A net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08806_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[19\]
+ net748 _04861_ _04875_ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__a211o_1
X_09786_ net349 _05330_ vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__nand2_1
XANTENNA__12456__A1 _03632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11259__A2 _07123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_134_Right_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08737_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[21\]
+ net666 net641 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout457_X net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08668_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[23\]
+ net796 net754 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout624_X net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08599_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[25\]
+ net592 _04669_ _04674_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[25\]
+ sky130_fd_sc_hd__o22a_2
XANTENNA__09710__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13005__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10630_ _06089_ _06635_ vssd1 vssd1 vccd1 vccd1 _06636_ sky130_fd_sc_hd__or2_1
XANTENNA__09624__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08326__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10561_ net382 _06570_ vssd1 vssd1 vccd1 vccd1 _06571_ sky130_fd_sc_hd__and2_1
XANTENNA__12844__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12300_ _03557_ _03575_ _03592_ vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__or3b_1
XFILLER_0_64_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13280_ net276 net2765 net434 vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10492_ _06467_ _06504_ net519 vssd1 vssd1 vccd1 vccd1 _06505_ sky130_fd_sc_hd__mux2_1
X_12231_ _08014_ _08018_ _03525_ vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_20_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10217__X _06243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08060__A1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[31\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12162_ _07920_ _07969_ _07962_ vssd1 vssd1 vccd1 vccd1 _07974_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11113_ _07079_ vssd1 vssd1 vccd1 vccd1 _07080_ sky130_fd_sc_hd__inv_2
XANTENNA__13675__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16970_ clknet_leaf_196_wb_clk_i _02600_ _00666_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_12093_ _07895_ _07903_ _07897_ vssd1 vssd1 vccd1 vccd1 _07905_ sky130_fd_sc_hd__a21oi_2
X_15921_ net1273 vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__inv_2
X_11044_ net964 _06691_ _07013_ vssd1 vssd1 vccd1 vccd1 _07014_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08899__B1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08363__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15852_ net1293 vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__inv_2
XANTENNA__09604__D net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14803_ net1216 vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__inv_2
XANTENNA__12447__A1 _03657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15783_ net1290 vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12995_ net562 _03698_ _03708_ vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__or3_4
X_17522_ clknet_leaf_113_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[25\]
+ _01218_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[25\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_99_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14734_ net1187 vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__inv_2
X_11946_ _07756_ _07757_ vssd1 vssd1 vccd1 vccd1 _07758_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17453_ clknet_leaf_49_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[21\]
+ _01149_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_14665_ net1222 vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__inv_2
X_11877_ _07652_ _07661_ _07688_ _07656_ vssd1 vssd1 vccd1 vccd1 _07689_ sky130_fd_sc_hd__a2bb2o_1
X_16404_ clknet_leaf_127_wb_clk_i _02034_ _00100_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_13616_ net2728 net296 net395 vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__mux2_1
X_17384_ clknet_leaf_49_wb_clk_i net1444 _01080_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10828_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[9\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06825_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09076__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14596_ net1227 vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__inv_2
XANTENNA__08236__C net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16335_ net1129 vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_45_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13547_ net2232 net292 net400 vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__mux2_1
XANTENNA__08823__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12754__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10759_ net1018 _04272_ _06051_ _06756_ vssd1 vssd1 vccd1 vccd1 _06757_ sky130_fd_sc_hd__a211o_1
XANTENNA__11511__X _07422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16266_ net1113 vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__inv_2
X_13478_ net275 net2661 net410 vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__mux2_1
X_18005_ clknet_leaf_82_wb_clk_i _03344_ _01701_ vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15217_ net1216 vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__inv_2
XFILLER_0_164_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12429_ _03605_ net1911 net215 vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__mux2_1
X_16197_ net1145 vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__inv_2
XANTENNA__12055__A team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[11\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15148_ net1077 vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__inv_2
XANTENNA__13585__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15079_ net1104 vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_71_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09000__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08354__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09640_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[1\]
+ net946 net930 net927 vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__and4_1
Xclkbuf_leaf_109_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_109_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_160_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09571_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[2\]
+ net944 net939 net936 vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__and4_1
XANTENNA__08106__A2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08522_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[26\]
+ net705 net604 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_69_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08453_ _04516_ _04519_ _04521_ _04531_ vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__or4_1
XFILLER_0_9_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14148__C net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08384_ _04458_ _04460_ _04462_ _04464_ vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__or4_1
XFILLER_0_163_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08814__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1061_A net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout417_A _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09005_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[14\]
+ net705 net641 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__a22o_1
XANTENNA__10184__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout205_X net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout786_A _04400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13495__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout510 net511 vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout521 net522 vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__buf_2
X_09907_ _05078_ _05101_ vssd1 vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__nand2_1
Xfanout532 _05633_ vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__clkbuf_2
Xfanout543 net545 vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__clkbuf_4
Xfanout554 net556 vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__clkbuf_4
Xfanout565 net567 vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__buf_2
Xfanout576 net577 vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__buf_2
X_09838_ _05863_ _05864_ _05866_ _05868_ vssd1 vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__or4_1
Xfanout598 net601 vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12839__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout741_X net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09769_ _05787_ _05790_ _05798_ _05799_ vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__or4_1
XANTENNA__17641__D team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout839_X net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11800_ _07580_ _07589_ _07593_ vssd1 vssd1 vccd1 vccd1 _07612_ sky130_fd_sc_hd__nand3_1
XANTENNA__09721__B net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12780_ net279 net2648 net488 vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__mux2_1
XANTENNA__08177__X _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09845__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11731_ _07538_ _07530_ _07519_ vssd1 vssd1 vccd1 vccd1 _07543_ sky130_fd_sc_hd__and3b_1
XFILLER_0_56_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11652__A2 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10359__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08337__B net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14450_ net1238 vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11662_ net31 net990 net917 net1801 vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__o22a_1
XFILLER_0_22_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09058__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13401_ net2025 net241 net419 vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__mux2_1
X_10613_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[9\] net906 net897
+ _06619_ vssd1 vssd1 vccd1 vccd1 _06620_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_64_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12574__S _03678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14381_ net1491 vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12601__A1 _07797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08805__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11593_ net2846 net1010 net345 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[31\]
+ vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16120_ net1134 vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10544_ net382 _06554_ vssd1 vssd1 vccd1 vccd1 _06555_ sky130_fd_sc_hd__and2_1
X_13332_ net219 net2746 net427 vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16051_ net1285 vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13263_ net199 net2820 net434 vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_31_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10475_ _06143_ _06145_ vssd1 vssd1 vccd1 vccd1 _06489_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15002_ net1058 vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__inv_2
X_12214_ _07476_ _07524_ _03508_ _07541_ vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__or4b_1
XANTENNA__09736__X _05768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13194_ net197 net2717 net352 vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_7_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08584__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12145_ _07955_ _07956_ vssd1 vssd1 vccd1 vccd1 _07957_ sky130_fd_sc_hd__nand2_1
XANTENNA__10391__A2 _06408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09184__A _05208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12076_ _07878_ _07882_ _07884_ _07886_ _07887_ vssd1 vssd1 vccd1 vccd1 _07888_ sky130_fd_sc_hd__o32ai_4
X_16953_ clknet_leaf_10_wb_clk_i _02583_ _00649_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09615__C net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11027_ _06999_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[7\] net568
+ vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__mux2_1
X_15904_ net1257 vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__inv_2
XANTENNA__10679__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16884_ clknet_leaf_128_wb_clk_i _02514_ _00580_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_202_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_202_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15835_ net1305 vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__inv_2
XANTENNA__12749__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15766_ net1297 vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__inv_2
XANTENNA__14290__B1 _05921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12978_ net269 net2209 net464 vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09836__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17505_ clknet_leaf_107_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[8\]
+ _01201_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_18367__1352 vssd1 vssd1 vccd1 vccd1 _18367__1352/HI net1352 sky130_fd_sc_hd__conb_1
X_14717_ net1087 vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11643__A2 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11929_ _07740_ vssd1 vssd1 vccd1 vccd1 _07741_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15697_ net1144 vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17436_ clknet_leaf_65_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[4\]
+ _01132_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_99_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09049__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14648_ net1200 vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14042__B1 _07451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_70_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_144_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12484__S net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17367_ clknet_leaf_42_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[31\]
+ _01063_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12337__X _03632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14579_ net1212 vssd1 vssd1 vccd1 vccd1 _00209_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16318_ net1138 vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17298_ clknet_leaf_125_wb_clk_i _02928_ _00994_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16249_ net1138 vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__clkbuf_4
XANTENNA_wire375_X net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__buf_2
Xoutput124 net124 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__buf_2
XFILLER_0_2_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09221__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10906__A1 _06214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput135 net135 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__buf_2
Xoutput146 net146 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
Xoutput157 net157 vssd1 vssd1 vccd1 vccd1 gpio_out[36] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08575__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput168 net168 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__clkbuf_4
Xoutput179 net179 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_110_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08327__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09623_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[2\]
+ net659 _05640_ _05645_ _05652_ vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout367_A net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09554_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[3\]
+ net710 net643 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[3\]
+ _05590_ vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__a221o_1
XANTENNA__09288__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10687__B _05949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09827__A2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08505_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[27\]
+ net816 net791 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09485_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[4\]
+ net819 net775 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[4\]
+ _05524_ vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__a221o_1
XFILLER_0_144_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1276_A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08436_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[28\]
+ net688 net678 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_77_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08367_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[30\]
+ net791 net775 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout701_A _04293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12595__A0 _03645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1064_X net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08298_ _04236_ _04240_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[21\]
+ _04151_ _04230_ vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__o2111a_1
XANTENNA__09460__B1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08173__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[10\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14336__A1 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14336__B2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10260_ _06159_ _06283_ net530 vssd1 vssd1 vccd1 vccd1 _06284_ sky130_fd_sc_hd__mux2_2
XANTENNA__09212__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout691_X net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout789_X net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08566__A2 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ net2390 net190 net541 vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__mux2_1
XANTENNA__09716__B net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_115_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11570__B2 _07438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1305 net1306 vssd1 vssd1 vccd1 vccd1 net1305 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout956_X net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout340 _03693_ vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__buf_2
XANTENNA__09515__A1 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout351 _03717_ vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__buf_4
Xfanout362 _05770_ vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__clkbuf_2
X_13950_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[3\] _03821_ _03822_
+ vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__nand3_1
Xfanout384 net387 vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__buf_8
XFILLER_0_89_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout395 _03732_ vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__buf_6
X_12901_ net240 net2131 net475 vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__mux2_1
X_13881_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[12\]
+ net560 net576 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[12\]
+ net987 vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__a221o_1
XANTENNA__12569__S net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10530__C1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15620_ net1171 vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__inv_2
X_12832_ net218 net2519 net482 vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__mux2_1
XANTENNA__09279__B1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09818__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15551_ net1117 vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12763_ net189 net2192 net489 vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14502_ net1208 vssd1 vssd1 vccd1 vccd1 _00132_ sky130_fd_sc_hd__inv_2
X_18270_ clknet_leaf_36_wb_clk_i _03499_ _01965_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[24\]
+ sky130_fd_sc_hd__dfrtp_4
X_11714_ _07522_ _07523_ _07525_ vssd1 vssd1 vccd1 vccd1 _07526_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15482_ net1147 vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__inv_2
XFILLER_0_167_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12694_ net193 net2965 net497 vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17221_ clknet_leaf_18_wb_clk_i _02851_ _00917_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_14433_ net1235 vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__inv_2
XANTENNA__13701__B _06743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11645_ net18 net991 net918 net1974 vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_42_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17152_ clknet_leaf_126_wb_clk_i _02782_ _00848_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput15 DAT_I[21] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14364_ _04083_ _04086_ _04090_ _04089_ _04088_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__o32a_1
X_11576_ net1949 net1004 net727 _07418_ vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__a22o_1
XANTENNA__12050__A2 _07468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput26 DAT_I[31] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_154_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09451__B1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput37 gpio_in[37] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_1
Xinput48 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_1
X_16103_ net1300 vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__inv_2
Xinput59 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13315_ net2578 net280 net428 vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__mux2_1
XANTENNA__14327__A1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10527_ _05833_ _05962_ _04279_ vssd1 vssd1 vccd1 vccd1 _06538_ sky130_fd_sc_hd__o21ai_1
X_17083_ clknet_leaf_193_wb_clk_i _02713_ _00779_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14327__B2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10118__A _05034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14295_ _04613_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[26\]
+ _04656_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[25\]
+ _04064_ vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_131_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16034_ net1282 vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__inv_2
XANTENNA__09907__A _05078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10458_ net334 _06309_ _06471_ _06472_ vssd1 vssd1 vccd1 vccd1 _06473_ sky130_fd_sc_hd__o211a_1
X_13246_ net270 net2906 net436 vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_90_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10389_ _05976_ _06406_ net889 vssd1 vssd1 vccd1 vccd1 _06407_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13177_ net270 net2445 net440 vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__mux2_1
XANTENNA__11561__B2 _07409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12128_ _07933_ _07937_ _07939_ vssd1 vssd1 vccd1 vccd1 _07940_ sky130_fd_sc_hd__or3_2
X_17985_ clknet_leaf_107_wb_clk_i _03324_ _01681_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_165_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12059_ net543 _07524_ _07867_ vssd1 vssd1 vccd1 vccd1 _07871_ sky130_fd_sc_hd__o21a_1
X_16936_ clknet_leaf_201_wb_clk_i _02566_ _00632_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12479__S net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16867_ clknet_leaf_199_wb_clk_i _02497_ _00563_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15818_ net1298 vssd1 vssd1 vccd1 vccd1 _01448_ sky130_fd_sc_hd__inv_2
X_16798_ clknet_leaf_185_wb_clk_i _02428_ _00494_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15749_ net1257 vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_138_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_193_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09270_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[9\]
+ net816 net788 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05320_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_103_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08221_ net883 net871 net867 vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__and3_1
X_17419_ clknet_leaf_50_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[19\]
+ _01115_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18399_ net915 vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_155_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12508__A _07840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08264__Y _04347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13103__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08152_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[4\] _04233_
+ vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__or2_4
XFILLER_0_99_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12041__A2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[20\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_151_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14318__A1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08083_ net1024 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__and2b_1
XANTENNA__08796__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14318__B2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[22\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12942__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_195_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_195_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08548__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_124_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_124_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08985_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[15\]
+ net814 net748 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[15\]
+ _05046_ vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout484_A _03703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12389__S net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout749_A net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08720__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09606_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[2\]
+ net885 net874 net860 vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__and4_1
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08168__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09537_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[3\]
+ net590 _05569_ _05574_ vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__o22ai_4
XANTENNA_fanout537_X net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1279_X net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08318__D net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09468_ _05508_ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08419_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[29\]
+ net828 net781 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout704_X net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12568__A0 _03605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09399_ _04350_ _05443_ _04246_ vssd1 vssd1 vccd1 vccd1 _05444_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_163_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13013__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11430_ team_05_WB.instance_to_wrap.wishbone.curr_state\[2\] team_05_WB.instance_to_wrap.wishbone.curr_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _07343_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09433__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11361_ _04216_ team_05_WB.instance_to_wrap.total_design.keypad0.next_rows\[3\] team_05_WB.instance_to_wrap.total_design.keypad0.next_rows\[2\]
+ vssd1 vssd1 vccd1 vccd1 _07302_ sky130_fd_sc_hd__and3_1
XANTENNA__11240__B1 _07124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08787__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12852__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13100_ net245 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[26\]
+ net451 vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__mux2_1
X_10312_ net531 _06235_ vssd1 vssd1 vccd1 vccd1 _06334_ sky130_fd_sc_hd__or2_1
X_14080_ _03946_ _03947_ _03931_ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__o21a_1
X_11292_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[1\] _07100_ _07126_
+ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[81\] _07251_ vssd1 vssd1
+ vccd1 vccd1 _07252_ sky130_fd_sc_hd__a221o_1
XANTENNA__08539__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10243_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[27\] _06101_ vssd1
+ vssd1 vccd1 vccd1 _06268_ sky130_fd_sc_hd__xor2_1
XFILLER_0_30_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13031_ net192 net2415 net456 vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__mux2_1
X_18366__1351 vssd1 vssd1 vccd1 vccd1 _18366__1351/HI net1351 sky130_fd_sc_hd__conb_1
XANTENNA__10346__A2 _06366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11543__B2 _07351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08944__C1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input45_A wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1102 net1103 vssd1 vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__buf_4
X_10174_ _06036_ _06045_ net521 vssd1 vssd1 vccd1 vccd1 _06201_ sky130_fd_sc_hd__mux2_1
Xfanout1113 net1120 vssd1 vssd1 vccd1 vccd1 net1113 sky130_fd_sc_hd__buf_4
Xfanout1124 net1126 vssd1 vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__buf_4
Xfanout1135 net1137 vssd1 vssd1 vccd1 vccd1 net1135 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13683__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1146 net1151 vssd1 vssd1 vccd1 vccd1 net1146 sky130_fd_sc_hd__buf_2
X_17770_ clknet_leaf_91_wb_clk_i _03113_ _01466_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1157 net1162 vssd1 vssd1 vccd1 vccd1 net1157 sky130_fd_sc_hd__buf_2
XANTENNA__12440__X _03671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14982_ net1208 vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__inv_2
Xfanout1168 net1170 vssd1 vssd1 vccd1 vccd1 net1168 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1179 net1181 vssd1 vssd1 vccd1 vccd1 net1179 sky130_fd_sc_hd__buf_4
X_16721_ clknet_leaf_118_wb_clk_i _02351_ _00417_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout192 _06217_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__clkbuf_2
X_13933_ _07451_ _03806_ _03807_ vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__and3_1
XFILLER_0_117_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08711__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16652_ clknet_leaf_2_wb_clk_i _02282_ _00348_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13864_ net1750 net982 _03768_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[3\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_53_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09612__D net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15603_ net1259 vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__inv_2
X_12815_ net279 net2269 net485 vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16583_ clknet_leaf_200_wb_clk_i _02213_ _00279_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13795_ net1595 net976 net725 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[6\]
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_83_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14808__A net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18322_ net1414 vssd1 vssd1 vccd1 vccd1 gpio_oeb[37] sky130_fd_sc_hd__buf_2
XANTENNA__13712__A net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15534_ net1132 vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08475__A1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12746_ net282 net2608 net492 vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18253_ clknet_leaf_38_wb_clk_i _03482_ _01948_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_38_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15465_ net1159 vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12328__A _07774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12677_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[12\]
+ net339 vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12559__A0 _03612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17204_ clknet_leaf_120_wb_clk_i _02834_ _00900_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14416_ net1092 vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__inv_2
X_18184_ clknet_leaf_39_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[5\]
+ _01879_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11628_ net1735 net1009 net344 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__a22o_1
X_15396_ net1227 vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__inv_2
XANTENNA__09424__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12047__B _07468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11589__D team_05_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11231__B1 _07128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08778__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17135_ clknet_leaf_137_wb_clk_i _02765_ _00831_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12762__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14347_ _04085_ _04090_ _04092_ _04119_ vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__or4_1
X_11559_ net1637 net1004 _07361_ net358 vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__a22o_1
Xhold607 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net2021 sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2032 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17066_ clknet_leaf_181_wb_clk_i _02696_ _00762_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold629 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net2043 sky130_fd_sc_hd__dlygate4sd3_1
X_14278_ net899 net921 _06907_ vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11378__S net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16017_ net1128 vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_59_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13229_ team_05_WB.instance_to_wrap.total_design.core.instr_fetch _04258_ _04262_
+ _03695_ vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__or4_4
XFILLER_0_97_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13593__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_6__f_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_6__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xhold1307 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 net2721 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12350__X _03645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08770_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[19\]
+ net699 net644 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[19\]
+ _04840_ vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__a221o_1
Xhold1318 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2732 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17968_ clknet_leaf_110_wb_clk_i _03307_ _01664_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__dfrtp_1
Xhold1329 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2743 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16919_ clknet_leaf_145_wb_clk_i _02549_ _00615_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_17899_ clknet_leaf_75_wb_clk_i _03242_ _01595_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08259__Y _04342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08702__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12937__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09322_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[8\]
+ net812 net784 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[8\]
+ _05364_ vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_122_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09663__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_153_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09253_ _05293_ _05300_ _05303_ vssd1 vssd1 vccd1 vccd1 _05304_ sky130_fd_sc_hd__or3_1
XFILLER_0_91_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout232_A _06367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08204_ _04232_ net962 _04271_ _04154_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__o311a_2
X_09184_ _05208_ _05235_ vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12014__A2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[23\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09415__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08135_ team_05_WB.instance_to_wrap.total_design.keypad0.key_counter\[3\] team_05_WB.instance_to_wrap.total_design.keypad0.key_counter\[2\]
+ team_05_WB.instance_to_wrap.total_design.keypad0.key_counter\[1\] team_05_WB.instance_to_wrap.total_design.keypad0.key_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__and4_1
XANTENNA__08154__C team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08769__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1141_A net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08066_ net1026 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[28\]
+ net971 _04182_ vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout699_A _04293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12722__A0 _06737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09194__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout487_X net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08941__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08968_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[15\]
+ net668 net629 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05031_ sky130_fd_sc_hd__a22o_1
XANTENNA__11289__B1 _07123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09282__A net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09713__C net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout654_X net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08899_ _04952_ _04960_ _04964_ net591 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[17\]
+ sky130_fd_sc_hd__o32a_4
XANTENNA__13008__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10930_ _06314_ _06768_ _06898_ _06920_ net565 vssd1 vssd1 vccd1 vccd1 _06921_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_92_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10500__A2 _06049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10861_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[10\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[10\]
+ _06857_ vssd1 vssd1 vccd1 vccd1 _06858_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout821_X net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12847__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_21_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_67_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12600_ net1658 _07798_ _03680_ vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13580_ net2872 net290 net396 vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__mux2_1
X_10792_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[24\] net1040 vssd1
+ vssd1 vccd1 vccd1 _06789_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10264__A1 _05577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12531_ _07798_ net1851 _03675_ vssd1 vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__mux2_1
XANTENNA__16616__Q team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15250_ net1238 vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__inv_2
X_12462_ net1874 _07798_ _03670_ vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09406__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14201_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[7\] _04003_
+ _04004_ vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__o21a_1
XANTENNA__13678__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11413_ net1891 _07326_ vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__xor2_1
XANTENNA__11213__B1 _07123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12582__S net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15181_ net1082 vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12393_ net1859 _03605_ net217 vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10567__A2 _06572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14132_ net2973 net504 net912 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[15\]
+ sky130_fd_sc_hd__and3_1
X_11344_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[13\] net509 net359
+ net979 vssd1 vssd1 vccd1 vccd1 _03396_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18307__1399 vssd1 vssd1 vccd1 vccd1 net1399 _18307__1399/LO sky130_fd_sc_hd__conb_1
X_14063_ team_05_WB.instance_to_wrap.CPU_DAT_O\[8\] net507 vssd1 vssd1 vccd1 vccd1
+ _03931_ sky130_fd_sc_hd__nand2_1
X_11275_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[42\] _07113_
+ _07116_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[74\] vssd1 vssd1
+ vccd1 vccd1 _07236_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09607__D _04296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_148_Right_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13014_ net283 net2325 net461 vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__mux2_1
XANTENNA__09185__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10226_ _05911_ _06249_ _06250_ vssd1 vssd1 vccd1 vccd1 _06251_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08393__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17822_ clknet_leaf_83_wb_clk_i _03165_ _01518_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[68\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13707__A net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08932__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10157_ net2156 net194 net540 vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold4 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[18\]
+ vssd1 vssd1 vccd1 vccd1 net1418 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_146_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17753_ clknet_leaf_98_wb_clk_i _03096_ _01449_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[63\]
+ sky130_fd_sc_hd__dfrtp_1
X_14965_ net1059 vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_85_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10088_ net515 _06115_ _06114_ vssd1 vssd1 vccd1 vccd1 _06116_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_59 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13916_ net1527 net981 _03794_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[29\]
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_50_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16704_ clknet_leaf_135_wb_clk_i _02334_ _00400_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_17684_ clknet_leaf_84_wb_clk_i _03027_ _01380_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[122\]
+ sky130_fd_sc_hd__dfrtp_1
X_14896_ net1183 vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16635_ clknet_leaf_193_wb_clk_i _02265_ _00331_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08239__C net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13847_ net1480 net580 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[25\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_18_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12757__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16566_ clknet_leaf_140_wb_clk_i _02196_ _00262_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13778_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[25\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[24\] team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[27\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[26\] vssd1
+ vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__or4_1
XFILLER_0_146_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15517_ net1147 vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_3_0_0_wb_clk_i_X clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18305_ net1397 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
XANTENNA__08999__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12729_ net194 net2616 net494 vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__mux2_1
X_16497_ clknet_leaf_123_wb_clk_i _02127_ _00193_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_18236_ clknet_leaf_57_wb_clk_i net1464 _01931_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15448_ net1168 vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13588__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18167_ clknet_leaf_46_wb_clk_i _03470_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.key_clk
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12492__S net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15379_ net1215 vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold404 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[124\] vssd1 vssd1
+ vccd1 vccd1 net1818 sky130_fd_sc_hd__dlygate4sd3_1
X_17118_ clknet_leaf_185_wb_clk_i _02748_ _00814_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold415 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[13\] vssd1 vssd1
+ vccd1 vccd1 net1829 sky130_fd_sc_hd__dlygate4sd3_1
X_18098_ clknet_leaf_54_wb_clk_i _03421_ _01794_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08271__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold426 net120 vssd1 vssd1 vccd1 vccd1 net1840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[10\] vssd1 vssd1
+ vccd1 vccd1 net1851 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold448 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[8\] vssd1
+ vssd1 vccd1 vccd1 net1862 sky130_fd_sc_hd__dlygate4sd3_1
Xhold459 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[117\] vssd1 vssd1
+ vccd1 vccd1 net1873 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17049_ clknet_leaf_15_wb_clk_i _02679_ _00745_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09940_ _05966_ _05968_ _05014_ vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout906 _04234_ vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09176__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout917 _07484_ vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__clkbuf_2
X_09871_ _04717_ _05899_ vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__nand2_1
Xfanout928 net929 vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_74_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout939 _04365_ vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__buf_2
X_08822_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[18\]
+ net606 net594 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[18\]
+ _04890_ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_146_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_146_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1104 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net2518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1115 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2529 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1126 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net2540 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10730__A2 _06729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1137 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2551 sky130_fd_sc_hd__dlygate4sd3_1
X_08753_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[21\]
+ net761 net734 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__a22o_1
Xhold1148 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net2562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1159 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2573 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_124_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10041__A net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08684_ net378 _04755_ vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__and2_1
XFILLER_0_136_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10494__A1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10976__A _04170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1091_A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18365__1350 vssd1 vssd1 vccd1 vccd1 _18365__1350/HI net1350 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_172_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11143__Y _07109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09305_ _04246_ _04348_ vssd1 vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__nor2_1
XANTENNA__09100__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11443__B1 _07348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout614_A _04318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09236_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[9\]
+ net653 net650 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13498__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09167_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[11\]
+ net833 net826 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[11\]
+ _05219_ vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout402_X net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14183__A team_05_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08118_ net1028 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[2\]
+ net972 _04208_ vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09098_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[12\]
+ net675 net632 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[12\]
+ _05154_ vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout983_A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09708__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08049_ net1043 vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1311_X net1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold960 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold971 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2385 sky130_fd_sc_hd__dlygate4sd3_1
X_11060_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[1\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[0\]
+ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[2\] vssd1 vssd1
+ vccd1 vccd1 _07027_ sky130_fd_sc_hd__and3_1
Xhold982 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 net2396 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09167__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold993 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 net2407 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout771_X net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout869_X net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10011_ _06036_ _06039_ net514 vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__mux2_1
XANTENNA__08914__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14750_ net1066 vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__inv_2
X_11962_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[0\] net993 vssd1
+ vssd1 vccd1 vccd1 _07774_ sky130_fd_sc_hd__nand2_4
XFILLER_0_99_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13701_ net900 _06743_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[1\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__10485__A1 _06494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10913_ _05908_ _05911_ vssd1 vssd1 vccd1 vccd1 _06906_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14681_ net1057 vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__inv_2
X_11893_ _07668_ _07704_ _07669_ vssd1 vssd1 vccd1 vccd1 _07705_ sky130_fd_sc_hd__o21a_1
XANTENNA__11481__S net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16420_ clknet_leaf_183_wb_clk_i _02050_ _00116_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13262__A team_05_WB.instance_to_wrap.total_design.core.instr_fetch vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13632_ net1958 net238 net391 vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__mux2_1
X_10844_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[0\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[0\]
+ _06839_ _06840_ vssd1 vssd1 vccd1 vccd1 _06841_ sky130_fd_sc_hd__and4_1
XFILLER_0_27_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16351_ clknet_leaf_156_wb_clk_i _01981_ _00047_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16346__Q team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13563_ net2204 net220 net399 vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10775_ team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.state\[0\] net1048
+ _06770_ team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.state\[1\] vssd1
+ vssd1 vccd1 vccd1 _06772_ sky130_fd_sc_hd__and4b_1
XFILLER_0_87_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15302_ net1280 vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12514_ _07789_ net1798 _03675_ vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__mux2_1
XANTENNA__09739__X _05770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16282_ net1255 vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13494_ net2182 net198 net405 vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__mux2_1
X_18021_ clknet_leaf_96_wb_clk_i _03360_ _01717_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15233_ net1224 vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__inv_2
X_12445_ net1757 _07789_ _03670_ vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13201__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15164_ net1074 vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__inv_2
X_12376_ net1896 _03646_ net217 vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__mux2_1
XANTENNA__09618__C net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14115_ net1687 net506 _03979_ vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__a21boi_2
X_11327_ net1920 net732 _07278_ _07285_ vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__o22a_1
X_15095_ net1101 vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__inv_2
X_14046_ _03888_ _03913_ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_157_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11258_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[11\] _07101_
+ _07128_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[67\] vssd1 vssd1
+ vccd1 vccd1 _07220_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10209_ _06158_ _06234_ net520 vssd1 vssd1 vccd1 vccd1 _06235_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11189_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[94\] _07096_
+ _07106_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[22\] vssd1 vssd1
+ vccd1 vccd1 _07154_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17805_ clknet_leaf_102_wb_clk_i _03148_ _01501_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[115\]
+ sky130_fd_sc_hd__dfrtp_1
X_15997_ net1128 vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10132__Y _06160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15652__A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17736_ clknet_leaf_94_wb_clk_i _03079_ _01432_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14948_ net1232 vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__inv_2
X_18330__1319 vssd1 vssd1 vccd1 vccd1 _18330__1319/HI net1319 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_141_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13662__A1 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_46 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12487__S net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17667_ clknet_leaf_90_wb_clk_i _03010_ _01363_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[105\]
+ sky130_fd_sc_hd__dfrtp_1
X_14879_ net1182 vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16618_ clknet_leaf_17_wb_clk_i _02248_ _00314_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_17598_ clknet_leaf_57_wb_clk_i _02969_ _01294_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08266__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[25\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13965__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16549_ clknet_leaf_179_wb_clk_i _02179_ _00245_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09021_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[14\]
+ net800 net750 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__a22o_1
X_18219_ clknet_leaf_80_wb_clk_i net1544 _01914_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13111__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09397__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold201 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[83\] vssd1 vssd1
+ vccd1 vccd1 net1615 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[112\] vssd1 vssd1
+ vccd1 vccd1 net1626 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold223 net96 vssd1 vssd1 vccd1 vccd1 net1637 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold234 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[0\] vssd1 vssd1
+ vccd1 vccd1 net1648 sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[73\] vssd1 vssd1
+ vccd1 vccd1 net1659 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12950__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold256 net148 vssd1 vssd1 vccd1 vccd1 net1670 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold267 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[17\] vssd1 vssd1
+ vccd1 vccd1 net1681 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold278 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[28\] vssd1 vssd1
+ vccd1 vccd1 net1692 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09923_ _05509_ _05950_ _05941_ vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_113_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09149__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold289 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[106\] vssd1 vssd1
+ vccd1 vccd1 net1703 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout703 _04292_ vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout714 _04288_ vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__buf_2
XANTENNA__08357__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17464__D net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout725 net726 vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_141_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout397_A _03731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout736 _04422_ vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__buf_4
XANTENNA__10323__X _06345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09854_ _05881_ _05882_ vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__nor2_1
Xfanout747 _04417_ vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__clkbuf_8
Xfanout758 net759 vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__buf_4
Xfanout769 net770 vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__clkbuf_8
X_08805_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[19\]
+ net794 net757 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__a22o_1
XANTENNA__11138__Y _07104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09785_ _05378_ _05815_ _05376_ vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_0_Left_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08736_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[21\]
+ net696 net612 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[21\]
+ _04807_ vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__a221o_1
XANTENNA__09321__A2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout731_A _07030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12397__S net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08667_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[23\]
+ net792 net772 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[23\]
+ _04737_ vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout352_X net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1094_X net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout829_A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18306__1398 vssd1 vssd1 vccd1 vccd1 net1398 _18306__1398/LO sky130_fd_sc_hd__conb_1
XFILLER_0_49_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08598_ _04661_ _04671_ _04672_ _04673_ vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__or4_1
XANTENNA__08176__A team_05_WB.instance_to_wrap.total_design.core.instr_fetch vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09710__D net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1261_X net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout617_X net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09559__X _05596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10560_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[12\] net906 _05736_
+ _06567_ _06569_ vssd1 vssd1 vccd1 vccd1 _06570_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_8_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17639__D team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09219_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[10\]
+ net768 net764 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[10\]
+ _05270_ vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09719__B net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08182__Y _04265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10491_ _06025_ _06038_ vssd1 vssd1 vccd1 vccd1 _06504_ sky130_fd_sc_hd__nand2_1
XANTENNA__12916__A0 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13021__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12230_ _08012_ _08018_ _08014_ vssd1 vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09388__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12392__A1 _07797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08596__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12161_ _07920_ _07969_ _07962_ vssd1 vssd1 vccd1 vccd1 _07973_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12860__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11112_ _07052_ _07058_ vssd1 vssd1 vccd1 vccd1 _07079_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_9_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12092_ _07903_ vssd1 vssd1 vccd1 vccd1 _07904_ sky130_fd_sc_hd__inv_2
Xhold790 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net2204 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08348__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15920_ net1265 vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__inv_2
X_11043_ net1046 _06703_ _07012_ net959 vssd1 vssd1 vccd1 vccd1 _07013_ sky130_fd_sc_hd__o211a_1
XANTENNA__10155__B1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15851_ net1306 vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__inv_2
X_14802_ net1238 vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15782_ net1272 vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__inv_2
XANTENNA__13644__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12994_ net307 net2102 net465 vssd1 vssd1 vccd1 vccd1 _02646_ sky130_fd_sc_hd__mux2_1
XANTENNA__10458__A1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1490 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2904 sky130_fd_sc_hd__dlygate4sd3_1
X_17521_ clknet_leaf_113_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[24\]
+ _01217_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[24\]
+ sky130_fd_sc_hd__dfrtp_4
X_14733_ net1082 vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__inv_2
XANTENNA__09312__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11945_ _07730_ _07738_ _07754_ _07734_ vssd1 vssd1 vccd1 vccd1 _07757_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_19_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08520__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17452_ clknet_leaf_50_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[20\]
+ _01148_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14664_ net1222 vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11876_ _07652_ _07662_ _07659_ vssd1 vssd1 vccd1 vccd1 _07688_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_60_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_28_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16403_ clknet_leaf_164_wb_clk_i _02033_ _00099_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13615_ net1994 net298 net395 vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__mux2_1
X_17383_ clknet_leaf_59_wb_clk_i net1433 _01079_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10827_ _06823_ vssd1 vssd1 vccd1 vccd1 _06824_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14595_ net1196 vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13720__A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16334_ net1126 vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13546_ net2019 net279 net400 vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10758_ _05802_ _06754_ vssd1 vssd1 vccd1 vccd1 _06756_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_109_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16265_ net1115 vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__inv_2
X_13477_ net273 net2312 net408 vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10689_ _05553_ _05807_ vssd1 vssd1 vccd1 vccd1 _06691_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_97_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18004_ clknet_leaf_82_wb_clk_i _03343_ _01700_ vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__dfrtp_1
X_15216_ net1093 vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__inv_2
X_12428_ net1623 _07797_ _03667_ vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09379__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16196_ net1145 vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11186__A2 _07119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12383__A1 _03632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12055__B _07379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08587__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15647__A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15147_ net1069 vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__inv_2
X_12359_ _03608_ _03631_ _03635_ _03637_ _03653_ vssd1 vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__o2111a_1
XANTENNA__12770__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15078_ net1209 vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_71_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14029_ _03892_ _03897_ vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_71_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09551__A2 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_160_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15382__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09570_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[2\]
+ net950 net939 net936 vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_160_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09839__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08521_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[26\]
+ net689 net658 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[26\]
+ _04595_ vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__a221o_1
X_17719_ clknet_leaf_76_wb_clk_i _03062_ _01415_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[93\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_149_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_149_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08511__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13106__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08452_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[28\]
+ net635 _04530_ net722 vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__a211o_1
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09067__A1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[25\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08383_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[30\]
+ net766 _04463_ net855 vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__a211o_1
XANTENNA__12945__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14726__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout312_A _06720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09004_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[14\]
+ net692 net646 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[14\]
+ _05063_ vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__a221o_1
XFILLER_0_143_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11177__A2 _07099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12374__A1 _03657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08578__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1221_A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_105_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_112_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout500 _07857_ vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout681_A _04301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout779_A net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout511 _06057_ vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__clkbuf_4
X_09906_ _05057_ _05058_ vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__nor2_2
Xfanout522 _05699_ vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__clkbuf_2
Xfanout544 net545 vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout1107_X net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout555 net556 vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__clkbuf_4
Xfanout566 net567 vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__buf_2
Xfanout577 _03764_ vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__buf_2
XANTENNA__09542__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09837_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[20\]
+ net814 net798 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[20\]
+ _05867_ vssd1 vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__a221o_1
Xfanout599 net601 vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout946_A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15292__A net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08750__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09768_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[0\]
+ net628 _05777_ _05780_ _05784_ vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_77_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08719_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[22\]
+ net789 net736 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout734_X net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09721__C net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09699_ _05731_ vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__inv_2
XANTENNA__08502__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13016__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11730_ net550 _07541_ vssd1 vssd1 vccd1 vccd1 _07542_ sky130_fd_sc_hd__nand2_2
XFILLER_0_95_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08337__C _04418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11661_ net32 net992 _07483_ net1693 vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__a22o_1
XANTENNA__12855__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13400_ net2967 net245 net419 vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__mux2_1
X_10612_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[9\] _06089_ vssd1
+ vssd1 vccd1 vccd1 _06619_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_25_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_54_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14380_ net1495 vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11592_ net994 _07472_ vssd1 vssd1 vccd1 vccd1 _07473_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_144_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_18_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13331_ net191 net2624 net426 vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10543_ _06549_ _06553_ vssd1 vssd1 vccd1 vccd1 _06554_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16050_ net1251 vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__inv_2
X_13262_ team_05_WB.instance_to_wrap.total_design.core.instr_fetch _04258_ _04262_
+ _03698_ vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__or4_4
X_10474_ net337 _06327_ _06333_ net334 _06487_ vssd1 vssd1 vccd1 vccd1 _06488_ sky130_fd_sc_hd__o221a_1
XFILLER_0_121_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11168__A2 _07102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15001_ net1058 vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08569__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12213_ _07523_ _08024_ vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__nand2_1
XANTENNA__13686__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09766__C1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12590__S net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13193_ net557 _04263_ vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__nand2_4
XFILLER_0_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_92_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09465__A net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12144_ _07944_ _07945_ _07951_ _07904_ vssd1 vssd1 vccd1 vccd1 _07956_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_124_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_63_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12075_ _07865_ _07868_ _07876_ vssd1 vssd1 vccd1 vccd1 _07887_ sky130_fd_sc_hd__and3_1
X_16952_ clknet_leaf_31_wb_clk_i _02582_ _00648_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09615__D net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11026_ net963 _06641_ _06998_ vssd1 vssd1 vccd1 vccd1 _06999_ sky130_fd_sc_hd__a21oi_1
X_15903_ net1294 vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__inv_2
XANTENNA__09533__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16883_ clknet_leaf_165_wb_clk_i _02513_ _00579_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13715__A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15834_ net1290 vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15765_ net1290 vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12977_ net261 net2582 net465 vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__mux2_1
XANTENNA__14290__A1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_183_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17504_ clknet_leaf_110_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[7\]
+ _01200_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11928_ _07730_ _07739_ vssd1 vssd1 vccd1 vccd1 _07740_ sky130_fd_sc_hd__nand2_1
X_14716_ net1095 vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15696_ net1144 vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_72_Left_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17435_ clknet_leaf_55_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[3\]
+ _01131_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_14647_ net1105 vssd1 vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12765__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11859_ _07670_ _07633_ _07634_ vssd1 vssd1 vccd1 vccd1 _07671_ sky130_fd_sc_hd__mux2_2
XFILLER_0_170_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17366_ clknet_leaf_35_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[30\]
+ _01062_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14578_ net1232 vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_136_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10603__A1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16317_ net1139 vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__inv_2
X_13529_ net2210 net191 net401 vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17297_ clknet_leaf_169_wb_clk_i _02927_ _00993_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16248_ net1133 vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13596__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__clkbuf_4
X_16179_ net1163 vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__inv_2
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__buf_2
XANTENNA__14281__A _06609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10367__B1 _05881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput125 net125 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__buf_2
XFILLER_0_10_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput136 net136 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__buf_2
Xoutput147 net147 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__clkbuf_4
XANTENNA__10906__A2 _06768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09375__A net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_81_Left_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput158 net158 vssd1 vssd1 vccd1 vccd1 gpio_out[37] sky130_fd_sc_hd__clkbuf_4
X_18305__1397 vssd1 vssd1 vccd1 vccd1 net1397 _18305__1397/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_110_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput169 net169 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__clkbuf_4
XANTENNA__09509__C1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08980__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14286__D_N _06387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09524__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire535_X net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08732__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09622_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[2\]
+ net652 _05639_ _05641_ _05646_ vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08278__X team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[21\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13608__A1 _06499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09553_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[3\]
+ net683 net594 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_108_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08504_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[27\]
+ net823 net765 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[27\]
+ _04581_ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_90_Left_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09484_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[4\]
+ net788 net765 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05524_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08435_ _04490_ _04511_ vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08366_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[30\]
+ net717 _04442_ _04446_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_92_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08799__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11151__Y _07117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08297_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[31\]
+ net851 net847 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[31\]
+ _04378_ vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08173__B team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14336__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_46_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_103_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout896_A net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14191__A _07031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1224_X net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10190_ _04265_ _06216_ vssd1 vssd1 vccd1 vccd1 _06217_ sky130_fd_sc_hd__and2_1
XANTENNA__09763__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout684_X net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09716__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1306 net1311 vssd1 vssd1 vccd1 vccd1 net1306 sky130_fd_sc_hd__buf_2
Xfanout330 _06705_ vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__clkbuf_2
Xfanout341 _03693_ vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__buf_4
Xfanout352 _03717_ vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__buf_6
XANTENNA__09515__A2 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout851_X net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout363 net364 vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__buf_2
XANTENNA__11322__A2 _07101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17652__D team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[19\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout385 net387 vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__buf_6
XANTENNA_fanout949_X net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout396 _03731_ vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__buf_6
X_12900_ net245 net2457 net475 vssd1 vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__mux2_1
XANTENNA__13094__X _03714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13880_ net1549 net983 _03776_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[11\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12831_ net189 net2534 net480 vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15550_ net1117 vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12762_ net195 net2908 net490 vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14501_ net1185 vssd1 vssd1 vccd1 vccd1 _00131_ sky130_fd_sc_hd__inv_2
X_11713_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[13\] net998 vssd1
+ vssd1 vccd1 vccd1 _07525_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15481_ net1158 vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12585__S net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12693_ net198 net2032 net497 vssd1 vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14366__A _04084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17220_ clknet_leaf_182_wb_clk_i _02850_ _00916_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_14432_ net1195 vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11644_ net19 net989 net916 net1725 vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_42_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12586__A1 _07793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17151_ clknet_leaf_151_wb_clk_i _02781_ _00847_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_3_5_0_wb_clk_i_X clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14363_ _04120_ _04135_ vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__or2_1
X_11575_ net1720 net1007 _07354_ _07453_ vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__a22o_1
XANTENNA__08254__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput16 DAT_I[22] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
Xinput27 DAT_I[3] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
X_16102_ net1130 vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput38 wb_rst_i vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_1
X_13314_ net2281 net283 net428 vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__mux2_1
Xinput49 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_1
X_17082_ clknet_leaf_12_wb_clk_i _02712_ _00778_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10526_ net2556 net276 net541 vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__mux2_1
XANTENNA__14327__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[5\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14294_ _04066_ vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16033_ net1251 vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_131_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13245_ net267 net2874 net436 vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10457_ _04970_ _06056_ _06298_ _06355_ vssd1 vssd1 vccd1 vccd1 _06472_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_90_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11010__A1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13176_ net269 net2215 net440 vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__mux2_1
X_10388_ _05883_ _05975_ vssd1 vssd1 vccd1 vccd1 _06406_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_1138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08962__B1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12127_ net547 _07657_ vssd1 vssd1 vccd1 vccd1 _07939_ sky130_fd_sc_hd__nand2_1
Xclkbuf_4_5__f_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_5__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_17984_ clknet_leaf_74_wb_clk_i _03323_ _01680_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09506__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12058_ net543 _07524_ vssd1 vssd1 vccd1 vccd1 _07870_ sky130_fd_sc_hd__nor2_1
X_16935_ clknet_leaf_201_wb_clk_i _02565_ _00631_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11313__A2 _07096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12510__A1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11009_ net1045 _06603_ _06984_ net959 vssd1 vssd1 vccd1 vccd1 _06985_ sky130_fd_sc_hd__o211a_1
XANTENNA__09642__B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16866_ clknet_leaf_8_wb_clk_i _02496_ _00562_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_15817_ net1277 vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16797_ clknet_leaf_111_wb_clk_i _02427_ _00493_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15748_ net1293 vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12495__S net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15679_ net1150 vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__inv_2
XANTENNA__08493__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08220_ net884 net862 net858 vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__and3_1
X_17418_ clknet_leaf_50_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[18\]
+ _01114_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_155_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18398_ net915 vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_155_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08151_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[4\] _04233_
+ vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__nor2_1
X_17349_ clknet_leaf_41_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[13\]
+ _01045_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08245__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12041__A3 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[21\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08082_ net1023 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[20\]
+ net970 _04190_ vssd1 vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__a22o_1
XANTENNA__14318__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[23\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12329__B2 _07774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08953__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08984_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[15\]
+ net822 net768 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1017_A _04347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12501__A1 _03666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11304__A2 _07110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout477_A net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_164_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_164_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_127_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09605_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[2\]
+ net877 net871 net857 vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__and4_1
XFILLER_0_79_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout644_A net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09536_ _05560_ _05570_ _05571_ _05573_ vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__or4_2
XANTENNA__11607__A3 _07472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13802__B net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09467_ _05506_ _05507_ vssd1 vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__nor2_2
XANTENNA__08484__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout811_A net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout432_X net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11162__X _07128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08418_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[29\]
+ net813 net774 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09398_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[26\] _04349_
+ vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__nand2_1
XFILLER_0_164_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08349_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[30\]
+ net706 net608 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10579__B1 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_128_Left_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11360_ _07290_ team_05_WB.instance_to_wrap.total_design.keypad0.next_rows\[2\] vssd1
+ vssd1 vccd1 vccd1 _07301_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17647__D team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[14\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout899_X net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10311_ _06227_ _06238_ net528 vssd1 vssd1 vccd1 vccd1 _06333_ sky130_fd_sc_hd__mux2_1
X_11291_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[9\] _07105_ _07127_
+ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[121\] vssd1 vssd1 vccd1
+ vccd1 _07251_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13030_ net195 net2363 net459 vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__mux2_1
XANTENNA__09197__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10242_ _06251_ _06265_ _06266_ _04275_ vssd1 vssd1 vccd1 vccd1 _06267_ sky130_fd_sc_hd__o31a_1
XFILLER_0_104_499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1103 net1107 vssd1 vssd1 vccd1 vccd1 net1103 sky130_fd_sc_hd__clkbuf_4
X_10173_ _06027_ _06039_ net519 vssd1 vssd1 vccd1 vccd1 _06200_ sky130_fd_sc_hd__mux2_1
Xfanout1114 net1120 vssd1 vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__buf_4
Xfanout1125 net1126 vssd1 vssd1 vccd1 vccd1 net1125 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1136 net1137 vssd1 vssd1 vccd1 vccd1 net1136 sky130_fd_sc_hd__buf_4
XANTENNA_input38_A wb_rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1147 net1150 vssd1 vssd1 vccd1 vccd1 net1147 sky130_fd_sc_hd__buf_4
Xfanout1158 net1161 vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__buf_4
X_14981_ net1203 vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__inv_2
XANTENNA__11484__S net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_137_Left_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1169 net1170 vssd1 vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_35_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16720_ clknet_leaf_124_wb_clk_i _02350_ _00416_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13932_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[4\] _03805_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__a21o_1
Xfanout193 _06184_ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13863_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[3\]
+ net560 net576 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[3\]
+ net987 vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__a221o_1
X_16651_ clknet_leaf_186_wb_clk_i _02281_ _00347_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15602_ net1258 vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__inv_2
X_12814_ net285 net2695 net485 vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__mux2_1
X_13794_ net1451 net975 net724 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[5\]
+ sky130_fd_sc_hd__and3_1
X_16582_ clknet_leaf_117_wb_clk_i _02212_ _00278_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09121__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18321_ net1413 vssd1 vssd1 vccd1 vccd1 gpio_oeb[36] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_83_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15533_ net1124 vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__inv_2
X_12745_ net276 net2811 net495 vssd1 vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__mux2_1
XANTENNA__08475__A2 _04552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18304__1396 vssd1 vssd1 vccd1 vccd1 net1396 _18304__1396/LO sky130_fd_sc_hd__conb_1
XFILLER_0_96_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13204__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15464_ net1159 vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__inv_2
X_18252_ clknet_leaf_39_wb_clk_i _03481_ _01947_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ net2969 net340 vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_146_Left_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17203_ clknet_leaf_168_wb_clk_i _02833_ _00899_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14415_ net1283 vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_133_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11627_ net2076 net1008 net345 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__a22o_1
X_18183_ clknet_leaf_41_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[4\]
+ _01878_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15395_ net1207 vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10129__A net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17134_ clknet_leaf_177_wb_clk_i _02764_ _00830_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_14346_ _04086_ _04087_ _04094_ _04095_ vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__or4_1
X_11558_ net727 _07452_ vssd1 vssd1 vccd1 vccd1 _07469_ sky130_fd_sc_hd__and2_1
XFILLER_0_163_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09956__A_N net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold608 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2022 sky130_fd_sc_hd__dlygate4sd3_1
Xwire583 net584 vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__clkbuf_1
X_10509_ _05104_ _05834_ vssd1 vssd1 vccd1 vccd1 _06521_ sky130_fd_sc_hd__xnor2_4
X_17065_ clknet_leaf_25_wb_clk_i _02695_ _00761_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14277_ _07025_ _07028_ _04051_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.lcd_en
+ sky130_fd_sc_hd__and3_1
Xhold619 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2033 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09637__B net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11489_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[22\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[22\]
+ net1031 vssd1 vssd1 vccd1 vccd1 _07400_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16016_ net1114 vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__inv_2
XANTENNA__09188__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13228_ _06766_ net2935 net351 vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__mux2_1
XANTENNA__09727__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08935__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13159_ net305 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[0\]
+ net444 vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__mux2_1
XANTENNA__10742__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_155_Left_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17967_ clknet_leaf_73_wb_clk_i _03306_ _01663_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__dfrtp_2
Xhold1308 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2722 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1319 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2733 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10151__X _06179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16918_ clknet_leaf_139_wb_clk_i _02548_ _00614_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08699__C1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17898_ clknet_leaf_95_wb_clk_i _03241_ _01594_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09360__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_0_wb_clk_i sky130_fd_sc_hd__clkbuf_16
X_16849_ clknet_leaf_123_wb_clk_i _02479_ _00545_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09112__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09321_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[8\]
+ net852 net740 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[8\]
+ _05358_ vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_122_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10738__S net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08466__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13114__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11470__A1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09252_ _05288_ _05289_ _05292_ _05302_ vssd1 vssd1 vccd1 vccd1 _05303_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_174_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12578__C_N _03659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08203_ net879 net875 net872 vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__nand3_4
XFILLER_0_172_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09183_ _05235_ vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__inv_2
XANTENNA__12953__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10039__A _04533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14734__A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_170_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08134_ team_05_WB.instance_to_wrap.total_design.keypad0.key_counter\[2\] _04220_
+ vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__and2_1
XFILLER_0_145_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08291__X _04373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10430__C1 _05924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08065_ net1025 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout1134_A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14172__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout594_A net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08967_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[15\]
+ net703 net594 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[15\]
+ _05029_ vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout761_A net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout382_X net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08898_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[17\]
+ net781 _04961_ _04963_ net854 vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09713__D net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout647_X net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10860_ _06822_ _06823_ _06856_ vssd1 vssd1 vccd1 vccd1 _06857_ sky130_fd_sc_hd__and3_1
X_09519_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[3\]
+ net806 net748 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05557_ sky130_fd_sc_hd__a22o_1
X_10791_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[24\] net1040 vssd1
+ vssd1 vccd1 vccd1 _06788_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout814_X net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08457__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13024__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12530_ net1694 _03604_ net208 vssd1 vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__mux2_1
XANTENNA__14347__C _04092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10264__A2 _06049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_61_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_81_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12461_ net1604 _03604_ net212 vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12863__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14200_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[7\] _04003_
+ net728 vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_124_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11412_ _07327_ _07336_ vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15180_ net1077 vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__inv_2
X_12392_ net1815 _07797_ _07852_ vssd1 vssd1 vccd1 vccd1 _03234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14131_ net1906 net502 net911 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[14\]
+ sky130_fd_sc_hd__and3_1
X_11343_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[14\] net509 net359
+ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[10\] vssd1 vssd1 vccd1
+ vccd1 _03397_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14062_ _03798_ _03930_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[7\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11274_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[122\] _07099_
+ _07108_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[90\] vssd1 vssd1
+ vccd1 vccd1 _07235_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08917__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13013_ net274 net2494 net463 vssd1 vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__mux2_1
X_10225_ _05911_ _06249_ _05924_ vssd1 vssd1 vccd1 vccd1 _06250_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_37_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17821_ clknet_leaf_100_wb_clk_i _03164_ _01517_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[67\]
+ sky130_fd_sc_hd__dfrtp_1
X_10156_ _04264_ _06183_ vssd1 vssd1 vccd1 vccd1 _06184_ sky130_fd_sc_hd__nor2_2
XANTENNA__11508__A _07414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold5 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[5\]
+ vssd1 vssd1 vccd1 vccd1 net1419 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17752_ clknet_leaf_93_wb_clk_i _03095_ _01448_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[62\]
+ sky130_fd_sc_hd__dfrtp_1
X_14964_ net1074 vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__inv_2
X_10087_ _06112_ _06113_ vssd1 vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_85_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09342__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16703_ clknet_leaf_155_wb_clk_i _02333_ _00399_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13915_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[29\]
+ net558 net574 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[29\]
+ net988 vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_50_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17683_ clknet_leaf_78_wb_clk_i _03026_ _01379_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08696__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14895_ net1240 vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload3_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13723__A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1086 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16634_ clknet_leaf_13_wb_clk_i _02264_ _00330_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13846_ net1472 net578 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[24\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_18_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13777_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[17\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[16\] team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[19\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[18\] vssd1
+ vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__or4_1
X_16565_ clknet_leaf_174_wb_clk_i _02195_ _00261_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08448__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10989_ net963 _06521_ net566 vssd1 vssd1 vccd1 vccd1 _06969_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_100_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18304_ net1396 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
X_15516_ net1144 vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12728_ net199 net2614 net494 vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__mux2_1
X_16496_ clknet_leaf_152_wb_clk_i _02126_ _00192_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18235_ clknet_leaf_57_wb_clk_i net1453 _01930_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15447_ net1168 vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__inv_2
XANTENNA__12773__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12659_ net2949 net341 vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__and2_1
XFILLER_0_170_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18166_ clknet_leaf_147_wb_clk_i _03469_ _01862_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15378_ net1240 vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17117_ clknet_leaf_111_wb_clk_i _02747_ _00813_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold405 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[35\] vssd1 vssd1
+ vccd1 vccd1 net1819 sky130_fd_sc_hd__dlygate4sd3_1
Xwire380 _04447_ vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__buf_4
X_14329_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[2\] net523
+ _04100_ _04101_ vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__a211o_1
Xhold416 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[77\] vssd1 vssd1
+ vccd1 vccd1 net1830 sky130_fd_sc_hd__dlygate4sd3_1
X_18097_ clknet_leaf_69_wb_clk_i _03420_ _01793_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[14\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08620__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08271__B net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold427 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1841 sky130_fd_sc_hd__dlygate4sd3_1
Xhold438 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[93\] vssd1 vssd1
+ vccd1 vccd1 net1852 sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[31\] vssd1 vssd1
+ vccd1 vccd1 net1863 sky130_fd_sc_hd__dlygate4sd3_1
X_17048_ clknet_leaf_30_wb_clk_i _02678_ _00744_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08908__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout907 _03994_ vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__clkbuf_4
X_09870_ _05888_ _05893_ _05898_ _05892_ _04757_ vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__a2111o_2
Xfanout918 _07483_ vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_74_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout929 _04376_ vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__buf_2
X_08821_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[18\]
+ net699 net668 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_146_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1105 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net2519 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1116 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net2530 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13109__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08752_ _04822_ _04823_ vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__nor2_1
Xhold1127 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2541 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10322__A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1138 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2552 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1149 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2563 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09333__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08683_ net378 _04755_ vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_124_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08687__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12948__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14729__A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08727__A _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09636__A1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout342_A _03693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08439__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09636__B2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09304_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[20\] net967
+ vssd1 vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout1084_A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09235_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[9\]
+ net630 net613 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09829__Y _05860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1251_A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout607_A _04320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09166_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[11\]
+ net794 net737 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08117_ net1028 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__and2b_1
X_09097_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[12\]
+ net710 net656 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08611__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_1__f_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1137_X net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09708__D net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08048_ net1 vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold950 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net2364 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout976_A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold961 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2375 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout597_X net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold972 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2386 sky130_fd_sc_hd__dlygate4sd3_1
Xhold983 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2397 sky130_fd_sc_hd__dlygate4sd3_1
Xhold994 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net2408 sky130_fd_sc_hd__dlygate4sd3_1
X_18303__1395 vssd1 vssd1 vccd1 vccd1 net1395 _18303__1395/LO sky130_fd_sc_hd__conb_1
X_10010_ _06037_ _06038_ vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout764_X net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09999_ _05123_ net365 vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__nand2_1
XANTENNA__13019__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09324__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11961_ net343 _07758_ _07772_ _07692_ _07750_ vssd1 vssd1 vccd1 vccd1 _07773_ sky130_fd_sc_hd__a32oi_4
XANTENNA__08678__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12858__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout931_X net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13700_ net899 _06756_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[0\]
+ sky130_fd_sc_hd__nor2_1
X_10912_ _06905_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[28\] net566
+ vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__mux2_1
X_14680_ net1210 vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__inv_2
XANTENNA__08196__X _04279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11892_ _07663_ _07665_ _07671_ vssd1 vssd1 vccd1 vccd1 _07704_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13631_ net2515 net244 net391 vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_50_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10843_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[1\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06840_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_80_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16350_ clknet_leaf_185_wb_clk_i _01980_ _00046_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13562_ net2006 net190 net398 vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__mux2_1
X_10774_ team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.state\[0\] team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06771_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_165_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08924__X _04989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12513_ net1692 _03651_ net209 vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__mux2_1
X_15301_ net1204 vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__inv_2
XANTENNA__13689__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16281_ net1255 vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__inv_2
XANTENNA__12593__S net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13493_ net557 _03694_ _03707_ vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__and3_1
XANTENNA__08850__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18020_ clknet_leaf_96_wb_clk_i _03359_ _01716_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12444_ net1713 _03651_ net213 vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15232_ net1196 vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11198__B1 _07109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15163_ net1100 vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__inv_2
X_12375_ net1707 _07793_ _07852_ vssd1 vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10945__B1 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14114_ _03978_ _03858_ _03977_ vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__or3b_1
XANTENNA__09618__D _04289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11326_ _07279_ _07281_ _07282_ _07284_ vssd1 vssd1 vccd1 vccd1 _07285_ sky130_fd_sc_hd__or4_1
XFILLER_0_120_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15094_ net1096 vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__inv_2
XANTENNA__13718__A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14045_ _03888_ _03913_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__and2b_1
X_11257_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[91\] _07096_
+ _07108_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[91\] _07218_
+ vssd1 vssd1 vccd1 vccd1 _07219_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_128_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09915__B _05801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10208_ _06171_ _06173_ vssd1 vssd1 vccd1 vccd1 _06234_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_52_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11188_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[14\] _07105_
+ _07126_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[86\] vssd1 vssd1
+ vccd1 vccd1 _07153_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_52_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17804_ clknet_leaf_77_wb_clk_i _03147_ _01500_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[114\]
+ sky130_fd_sc_hd__dfrtp_1
X_10139_ net379 net368 vssd1 vssd1 vccd1 vccd1 _06167_ sky130_fd_sc_hd__nand2_1
X_15996_ net1129 vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__inv_2
XANTENNA__09315__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17735_ clknet_leaf_86_wb_clk_i _03078_ _01431_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12768__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14947_ net1208 vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__inv_2
XANTENNA__08669__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17570__D team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09650__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17666_ clknet_leaf_98_wb_clk_i _03009_ _01362_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[104\]
+ sky130_fd_sc_hd__dfrtp_1
X_14878_ net1074 vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16617_ clknet_leaf_20_wb_clk_i _02247_ _00313_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13829_ net1933 net582 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[7\]
+ sky130_fd_sc_hd__and2_1
X_17597_ clknet_leaf_56_wb_clk_i _02968_ _01293_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12622__A0 _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16548_ clknet_leaf_183_wb_clk_i _02178_ _00244_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09094__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13599__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14284__A _06481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12356__X _03651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16479_ clknet_leaf_155_wb_clk_i _02109_ _00175_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08841__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09020_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[26\] net967
+ net955 _05080_ _04345_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[14\]
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_54_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18218_ clknet_leaf_79_wb_clk_i net1531 _01913_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11189__B1 _07106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18149_ clknet_leaf_116_wb_clk_i _03452_ _01845_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold202 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[95\] vssd1 vssd1
+ vccd1 vccd1 net1616 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_117_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09251__C1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold213 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[15\] vssd1 vssd1
+ vccd1 vccd1 net1627 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold224 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[0\] vssd1 vssd1
+ vccd1 vccd1 net1638 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09665__X team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold235 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[86\] vssd1 vssd1
+ vccd1 vccd1 net1649 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold246 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[113\] vssd1 vssd1
+ vccd1 vccd1 net1660 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_148_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold257 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[7\] vssd1 vssd1
+ vccd1 vccd1 net1671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 net127 vssd1 vssd1 vccd1 vccd1 net1682 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold279 team_05_WB.instance_to_wrap.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 net1693
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ _05509_ _05950_ vssd1 vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout704 _04292_ vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__buf_2
Xfanout715 _04286_ vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__buf_8
Xfanout726 _03759_ vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09554__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_165_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09853_ net360 _05879_ vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__and2_1
Xfanout737 net738 vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_165_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout748 net751 vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__buf_6
Xfanout759 _04412_ vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__buf_4
X_08804_ _04867_ _04869_ _04871_ _04873_ vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__or4_1
X_09784_ _05422_ _05814_ _05420_ vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__a21o_1
X_08735_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[21\]
+ net657 net634 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10987__A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11435__X _07348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1299_A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08666_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[23\]
+ net831 net812 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__a22o_1
XANTENNA__09560__B _05596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11154__Y _07120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08597_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[25\]
+ net851 net848 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[25\]
+ _04660_ vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout724_A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12613__A0 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_134_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_9_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13302__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09218_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[10\]
+ net814 net794 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10490_ net369 _06062_ vssd1 vssd1 vccd1 vccd1 _06503_ sky130_fd_sc_hd__nand2_2
XANTENNA__09719__C net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_101_Left_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09149_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[11\]
+ net676 net625 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[11\]
+ _05193_ vssd1 vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_20_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1030 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12160_ _07927_ _07929_ _07971_ vssd1 vssd1 vccd1 vccd1 _07972_ sky130_fd_sc_hd__nand3_1
XFILLER_0_130_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11111_ _07063_ _07067_ vssd1 vssd1 vccd1 vccd1 _07078_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_9_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12091_ _07893_ _07898_ _07900_ vssd1 vssd1 vccd1 vccd1 _07903_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_9_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold780 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2194 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13877__C1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold791 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 net2205 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09545__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11042_ _06834_ _06847_ _06848_ _07011_ vssd1 vssd1 vccd1 vccd1 _07012_ sky130_fd_sc_hd__a31o_1
XANTENNA__10155__A1 _04176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10155__B2 _06179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13892__A2 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15850_ net1298 vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_110_Left_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input20_A DAT_I[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14801_ net1192 vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__inv_2
XANTENNA__12588__S net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15781_ net1256 vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__inv_2
X_12993_ net326 net2310 net464 vssd1 vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11492__S net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17520_ clknet_leaf_72_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[23\]
+ _01216_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1480 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2894 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1491 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2905 sky130_fd_sc_hd__dlygate4sd3_1
X_14732_ net1071 vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__inv_2
X_11944_ _07752_ _07754_ _07755_ vssd1 vssd1 vccd1 vccd1 _07756_ sky130_fd_sc_hd__or3_2
XANTENNA_clkbuf_leaf_173_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_54_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11064__Y _07031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17451_ clknet_leaf_50_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[19\]
+ _01147_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11875_ _07685_ _07686_ vssd1 vssd1 vccd1 vccd1 _07687_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14663_ net1105 vssd1 vssd1 vccd1 vccd1 _00293_ sky130_fd_sc_hd__inv_2
XANTENNA_output107_A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16402_ clknet_leaf_123_wb_clk_i _02032_ _00098_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12604__A0 _03666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10826_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[10\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06823_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13614_ net2081 net287 net392 vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__mux2_1
X_17382_ clknet_leaf_60_wb_clk_i net1441 _01078_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14594_ net1204 vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__inv_2
XANTENNA__09076__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13720__B _06408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16333_ net1113 vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__inv_2
X_13545_ net2169 net284 net401 vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__mux2_1
XANTENNA__08284__B1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10757_ _04158_ _05802_ _06051_ _06754_ vssd1 vssd1 vccd1 vccd1 _06755_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_45_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08823__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13212__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16264_ net1113 vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__inv_2
X_13476_ net267 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[16\]
+ net408 vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10688_ net890 _06689_ vssd1 vssd1 vccd1 vccd1 _06690_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_97_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12336__B _07475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18003_ clknet_leaf_82_wb_clk_i _03342_ _01699_ vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12427_ net1729 _07798_ _03667_ vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__mux2_1
X_15215_ net1281 vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__inv_2
X_16195_ net1145 vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10137__A _04656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12055__C _07465_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12358_ _03638_ _03639_ _03640_ _03652_ vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__o31a_1
XFILLER_0_2_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15146_ net1121 vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10154__A1_N team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[30\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17565__D team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11309_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[72\] _07109_
+ _07130_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[96\] vssd1 vssd1
+ vccd1 vccd1 _07268_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15077_ net1184 vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__inv_2
XANTENNA__09645__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12289_ _08008_ _03583_ vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__nor2_1
X_14028_ _03892_ _03897_ vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_71_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_0__f_wb_clk_i_X clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09000__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10697__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_160_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12498__S _03673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14279__A _06706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15979_ net1304 vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08520_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[26\]
+ net667 net662 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[26\]
+ _04596_ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__a221o_1
X_17718_ clknet_leaf_78_wb_clk_i _03061_ _01414_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[92\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_69_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08451_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[28\]
+ net702 net639 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__a22o_1
X_17649_ clknet_leaf_54_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[16\]
+ _01345_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08382_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[30\]
+ net796 net762 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_189_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_189_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_45_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18302__1394 vssd1 vssd1 vccd1 vccd1 net1394 _18302__1394/LO sky130_fd_sc_hd__conb_1
XFILLER_0_46_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08814__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13122__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_118_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_118_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09003_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[14\]
+ net662 net612 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_115_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12961__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout305_A net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11031__C1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10334__X _06355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout501 _07515_ vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09527__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11149__Y _07115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout512 net515 vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__clkbuf_4
X_09905_ _04989_ _05011_ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__and2_1
Xfanout545 net546 vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout674_A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout556 _05925_ vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__clkbuf_4
Xfanout567 _06774_ vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__dlymetal6s2s_1
X_09836_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[20\]
+ net810 net741 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1002_X net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout578 net580 vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__clkbuf_2
XANTENNA__17561__Q team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout462_X net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout841_A net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09767_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[0\]
+ net607 _05773_ _05782_ _05785_ vssd1 vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__a2111o_1
X_08718_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[22\]
+ net773 net757 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[22\]
+ _04790_ vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__a221o_1
XFILLER_0_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09698_ _05725_ _05727_ _05730_ net716 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__o32a_4
XFILLER_0_96_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09721__D net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08649_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[23\]
+ net713 net697 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__a22o_1
X_11660_ net33 net990 net917 net1731 vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__o22a_1
XANTENNA__09058__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10611_ _06610_ _06616_ _06617_ net537 vssd1 vssd1 vccd1 vccd1 _06618_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_25_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12062__A1 _07478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11591_ team_05_WB.instance_to_wrap.wishbone.curr_state\[2\] _07452_ _07471_ vssd1
+ vssd1 vccd1 vccd1 _07472_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_25_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08805__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13032__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13330_ net193 net2111 net426 vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__mux2_1
XANTENNA__14339__B1 _05165_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10542_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[13\] net906 net968
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[13\] _06552_ vssd1
+ vssd1 vccd1 vccd1 _06553_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13261_ net308 net2278 net436 vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__mux2_1
XANTENNA__12871__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10473_ _05015_ net511 _06324_ _06355_ _06486_ vssd1 vssd1 vccd1 vccd1 _06487_ sky130_fd_sc_hd__o221a_1
XFILLER_0_134_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15000_ net1200 vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__inv_2
X_12212_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[14\] team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[6\]
+ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[5\] team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[4\]
+ vssd1 vssd1 vccd1 vccd1 _08024_ sky130_fd_sc_hd__and4b_1
XFILLER_0_32_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13192_ net307 net2612 net440 vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__mux2_1
XANTENNA_input68_A wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11487__S _07345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12143_ _07903_ _07948_ vssd1 vssd1 vccd1 vccd1 _07955_ sky130_fd_sc_hd__or2_1
Xclkbuf_4_4__f_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_4__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__13314__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12074_ _07865_ _07877_ _07876_ vssd1 vssd1 vccd1 vccd1 _07886_ sky130_fd_sc_hd__a21oi_2
X_16951_ clknet_leaf_143_wb_clk_i _02581_ _00647_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15902_ net1267 vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__inv_2
X_11025_ net1045 _06653_ _06997_ net959 vssd1 vssd1 vccd1 vccd1 _06998_ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10679__A2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16882_ clknet_leaf_126_wb_clk_i _02512_ _00578_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15833_ net1295 vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__inv_2
XANTENNA__13715__B _06500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17471__Q team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13207__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15764_ net1300 vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11628__B2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12976_ net265 net2537 net465 vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14290__A2 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17503_ clknet_leaf_114_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[6\]
+ _01199_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_14715_ net1098 vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__inv_2
X_11927_ _07731_ _07732_ _07734_ _07736_ vssd1 vssd1 vccd1 vccd1 _07739_ sky130_fd_sc_hd__a22o_1
X_15695_ net1144 vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13731__A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17434_ clknet_leaf_69_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[2\]
+ _01130_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14646_ net1084 vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__inv_2
XANTENNA__09049__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11858_ _07619_ _07633_ vssd1 vssd1 vccd1 vccd1 _07670_ sky130_fd_sc_hd__nand2_1
XANTENNA__14042__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10809_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[16\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06806_ sky130_fd_sc_hd__nand2_1
X_17365_ clknet_leaf_37_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[29\]
+ _01061_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08257__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11789_ _07600_ vssd1 vssd1 vccd1 vccd1 _07601_ sky130_fd_sc_hd__inv_2
X_14577_ net1188 vssd1 vssd1 vccd1 vccd1 _00207_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_136_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16316_ net1125 vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10603__A2 _06609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13528_ net2213 net195 net402 vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__mux2_1
X_17296_ clknet_leaf_124_wb_clk_i _02926_ _00992_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16247_ net1132 vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12781__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13459_ net2721 net305 net412 vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__clkbuf_4
X_16178_ net1163 vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__inv_2
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__buf_2
XANTENNA__14281__B _06623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09221__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput126 net126 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__clkbuf_4
Xoutput137 net137 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__buf_2
Xoutput148 net148 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__clkbuf_4
X_15129_ net1051 vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_110_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput159 net159 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_110_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_162_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13069__A0 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09621_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[2\]
+ net621 net607 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__a22o_1
XANTENNA__13117__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09552_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[3\]
+ net675 net668 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[3\]
+ _05579_ vssd1 vssd1 vccd1 vccd1 _05589_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10330__A net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11619__B2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[11\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09288__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08503_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[27\]
+ net796 net779 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__a22o_1
X_09483_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[4\]
+ net842 net791 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[4\]
+ _05522_ vssd1 vssd1 vccd1 vccd1 _05523_ sky130_fd_sc_hd__a221o_1
XANTENNA__08496__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12956__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout255_A _06442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08434_ _04512_ vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11432__Y _07345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08248__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08365_ _04432_ _04433_ _04444_ _04445_ vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__or4_1
XFILLER_0_163_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10329__X _06350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout422_A net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14175__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10055__B1 _04275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08296_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[31\]
+ net842 net838 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__a22o_1
XANTENNA__09460__A2 _04366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout210_X net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout308_X net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09212__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout791_A net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout889_A _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08420__B1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_86_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_30_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09716__D net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1307 net1309 vssd1 vssd1 vccd1 vccd1 net1307 sky130_fd_sc_hd__buf_4
Xfanout320 _06671_ vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11307__B1 _07129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout677_X net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_15_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout331 _06705_ vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__buf_1
Xfanout342 _03693_ vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__clkbuf_4
Xfanout353 _03717_ vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__buf_2
Xfanout364 _05770_ vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__buf_2
Xfanout386 net387 vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__clkbuf_8
X_09819_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[20\]
+ net703 net695 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[20\]
+ _05843_ vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__a221o_1
Xfanout397 _03731_ vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10530__A1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout844_X net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13027__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12830_ net194 net2345 net481 vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12761_ net199 net2447 net490 vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__mux2_1
XANTENNA__12866__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08487__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14500_ net1228 vssd1 vssd1 vccd1 vccd1 _00130_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11712_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[13\] net998 vssd1
+ vssd1 vccd1 vccd1 _07524_ sky130_fd_sc_hd__and2_1
X_15480_ net1158 vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__inv_2
X_12692_ _04262_ net563 _03695_ vssd1 vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__or3_1
XANTENNA__14366__B _04091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11643_ net20 net991 net918 net1936 vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__a22o_1
X_14431_ net1178 vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_42_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17150_ clknet_leaf_184_wb_clk_i _02780_ _00846_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11574_ net920 _07354_ _07427_ net1007 net1591 vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__a32o_1
X_14362_ _04093_ _04110_ _04121_ _04134_ vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__o22a_1
XANTENNA__09451__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput17 DAT_I[23] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
X_16101_ net1309 vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__inv_2
Xinput28 DAT_I[4] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
Xinput39 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
X_13313_ net2514 net276 net430 vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10525_ _04265_ _06536_ vssd1 vssd1 vccd1 vccd1 _06537_ sky130_fd_sc_hd__and2_1
X_17081_ clknet_leaf_6_wb_clk_i _02711_ _00777_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14293_ _04573_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13244_ net261 net2356 net437 vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__mux2_1
XANTENNA__09739__B1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16032_ net1287 vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_131_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10456_ net1018 _04968_ _04969_ net551 vssd1 vssd1 vccd1 vccd1 _06471_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_131_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09203__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11546__B1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11010__A2 _06591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13175_ net261 net2903 net440 vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__mux2_1
X_10387_ net2080 net247 net540 vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__mux2_1
X_12126_ net544 _07658_ vssd1 vssd1 vccd1 vccd1 _07938_ sky130_fd_sc_hd__nor2_1
X_17983_ clknet_leaf_107_wb_clk_i _03322_ _01679_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__dfrtp_1
XANTENNA__13726__A net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12057_ _07868_ vssd1 vssd1 vccd1 vccd1 _07869_ sky130_fd_sc_hd__inv_2
X_16934_ clknet_leaf_117_wb_clk_i _02564_ _00630_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_18301__1393 vssd1 vssd1 vccd1 vccd1 net1393 _18301__1393/LO sky130_fd_sc_hd__conb_1
XFILLER_0_165_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11008_ _04170_ _06857_ _06983_ vssd1 vssd1 vccd1 vccd1 _06984_ sky130_fd_sc_hd__or3b_1
X_16865_ clknet_leaf_148_wb_clk_i _02495_ _00561_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09642__C net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15816_ net1276 vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__inv_2
X_16796_ clknet_leaf_158_wb_clk_i _02426_ _00492_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15747_ net1301 vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_29_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08478__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12776__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12959_ net322 net2750 net471 vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_138_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15678_ net1154 vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09690__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17417_ clknet_leaf_50_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[17\]
+ _01113_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14629_ net1184 vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__inv_2
XANTENNA__10296__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18397_ net1371 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_155_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_155_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10037__B1 _06060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08150_ net1022 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[5\]
+ _04231_ vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__or3_4
XFILLER_0_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17348_ clknet_leaf_39_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[12\]
+ _01044_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12041__A4 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[24\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08081_ net1023 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[20\]
+ vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__and2b_1
XFILLER_0_67_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12364__X _03659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17279_ clknet_leaf_156_wb_clk_i _02909_ _00975_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08650__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14292__A _04613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_wire380_X net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13400__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_0_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08402__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08983_ _05039_ _05041_ _05042_ _05044_ vssd1 vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__or4_1
XANTENNA__10760__A1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_127_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09604_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[2\]
+ net885 net869 net864 vssd1 vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_127_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09535_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[3\]
+ net802 net764 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[3\]
+ _05572_ vssd1 vssd1 vccd1 vccd1 _05573_ sky130_fd_sc_hd__a221o_1
XANTENNA__08469__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1281_A net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09130__A1 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_133_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_133_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout637_A _04312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09466_ net374 _05505_ vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_947 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13802__C net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08417_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[29\]
+ net808 net797 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__a22o_1
X_09397_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[6\]
+ net715 _05436_ _05441_ vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_136_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout804_A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout425_X net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08184__B net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08348_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[30\]
+ net692 net684 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__a22o_1
XANTENNA__09848__X team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[20\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09433__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11240__A2 _07110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08279_ net573 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[21\] vssd1
+ vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__nor2_1
XFILLER_0_144_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10310_ _04717_ net552 _06055_ _05898_ _06331_ vssd1 vssd1 vccd1 vccd1 _06332_ sky130_fd_sc_hd__o221a_1
XANTENNA__13310__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11290_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[17\] _07106_
+ _07128_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[65\] vssd1 vssd1
+ vccd1 vccd1 _07250_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout794_X net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10241_ _06049_ _06257_ _06258_ _05910_ vssd1 vssd1 vccd1 vccd1 _06266_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__18402__A net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10172_ _06198_ vssd1 vssd1 vccd1 vccd1 _06199_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout961_X net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1104 net1106 vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__buf_4
XANTENNA__10751__A1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1115 net1120 vssd1 vssd1 vccd1 vccd1 net1115 sky130_fd_sc_hd__buf_2
Xfanout1126 net1127 vssd1 vssd1 vccd1 vccd1 net1126 sky130_fd_sc_hd__clkbuf_2
Xfanout1137 net1177 vssd1 vssd1 vccd1 vccd1 net1137 sky130_fd_sc_hd__clkbuf_2
X_14980_ net1236 vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__inv_2
Xfanout1148 net1150 vssd1 vssd1 vccd1 vccd1 net1148 sky130_fd_sc_hd__buf_2
Xfanout1159 net1160 vssd1 vssd1 vccd1 vccd1 net1159 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13931_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[4\] team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[1\]
+ _03805_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__nand3_1
Xfanout194 _06184_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__dlymetal6s2s_1
X_16650_ clknet_leaf_17_wb_clk_i _02280_ _00346_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13862_ net1808 net982 _03767_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[2\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_87_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15601_ net1253 vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__inv_2
X_12813_ net276 net2617 net486 vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__mux2_1
XANTENNA__12596__S _03680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16581_ clknet_leaf_175_wb_clk_i _02211_ _00277_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13793_ net1571 net976 net725 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[4\]
+ sky130_fd_sc_hd__and3_1
X_18320_ net1412 vssd1 vssd1 vccd1 vccd1 gpio_oeb[35] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_83_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15532_ net1139 vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ net272 net2757 net492 vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18251_ clknet_leaf_38_wb_clk_i _03480_ _01946_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13205__A0 _06422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15463_ net1160 vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[14\]
+ net342 vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__and2_1
XFILLER_0_166_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17202_ clknet_leaf_133_wb_clk_i _02832_ _00898_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_14414_ net1191 vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18182_ clknet_leaf_42_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[3\]
+ _01877_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11626_ net2507 net1008 net344 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_133_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15394_ net1226 vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09424__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10129__B net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17133_ clknet_leaf_160_wb_clk_i _02763_ _00829_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11231__A2 _07104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14345_ _04099_ _04111_ _04116_ _04117_ vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__nand4_1
X_11557_ _07389_ _07458_ _07462_ _07464_ vssd1 vssd1 vccd1 vccd1 _07468_ sky130_fd_sc_hd__or4_4
XFILLER_0_135_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08632__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13220__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10508_ net888 _06519_ vssd1 vssd1 vccd1 vccd1 _06520_ sky130_fd_sc_hd__nor2_1
X_17064_ clknet_leaf_204_wb_clk_i _02694_ _00760_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold609 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net2023 sky130_fd_sc_hd__dlygate4sd3_1
Xwire584 _05763_ vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__clkbuf_1
X_14276_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[3\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[2\]
+ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[4\] vssd1 vssd1
+ vccd1 vccd1 _04051_ sky130_fd_sc_hd__a21oi_1
X_11488_ _07396_ _07392_ _07394_ _07398_ vssd1 vssd1 vccd1 vccd1 _07399_ sky130_fd_sc_hd__nand4b_1
XFILLER_0_150_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09637__C net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16015_ net1112 vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__inv_2
X_10439_ net337 _06278_ _06280_ net334 _06454_ vssd1 vssd1 vccd1 vccd1 _06455_ sky130_fd_sc_hd__o221a_1
X_13227_ net327 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[1\]
+ net351 vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10145__A _04533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09593__D1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13158_ net325 net1962 net444 vssd1 vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__mux2_1
X_12109_ _07466_ _07600_ _07919_ _07913_ _07912_ vssd1 vssd1 vccd1 vccd1 _07921_ sky130_fd_sc_hd__a32o_1
X_17966_ clknet_leaf_106_wb_clk_i _03305_ _01662_ vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__dfrtp_1
X_13089_ net331 net2221 net454 vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__mux2_1
Xhold1309 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net2723 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16917_ clknet_leaf_23_wb_clk_i _02547_ _00613_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11298__A2 _07118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12495__A1 _03664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17897_ clknet_leaf_105_wb_clk_i _03240_ _01593_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16848_ clknet_leaf_137_wb_clk_i _02478_ _00544_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_105_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16779_ clknet_leaf_187_wb_clk_i _02409_ _00475_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14287__A _06350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09320_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[8\]
+ net789 net735 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[8\]
+ _05356_ vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09663__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09251_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[9\]
+ net674 _05301_ net721 vssd1 vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__a211o_1
XFILLER_0_8_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11470__A2 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08871__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08202_ net879 net874 net871 vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__and3_4
XFILLER_0_90_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09182_ net570 net535 _05215_ vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09415__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_170_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08133_ team_05_WB.instance_to_wrap.total_design.keypad0.key_counter\[1\] team_05_WB.instance_to_wrap.total_design.keypad0.key_counter\[0\]
+ _04219_ vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11222__A2 _07120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08623__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout218_A net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13130__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08064_ net1025 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[29\]
+ net971 _04181_ vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1127_A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11438__X _07351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08966_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[15\]
+ net672 net656 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__a22o_1
XANTENNA__11157__Y _07123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12486__A1 _03610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11289__A2 _07099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout754_A net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08897_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[17\]
+ net815 net790 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[17\]
+ _04962_ vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_162_Right_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_40_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout921_A _05213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout542_X net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13305__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09518_ _05556_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[3\]
+ sky130_fd_sc_hd__inv_2
X_10790_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[25\] net1040 vssd1
+ vssd1 vccd1 vccd1 _06787_ sky130_fd_sc_hd__and2_1
XANTENNA__09654__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09449_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[5\]
+ net776 net766 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__a22o_1
XANTENNA__08862__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout807_X net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12460_ net1785 _03664_ net213 vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__mux2_1
XANTENNA__09406__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18300__1392 vssd1 vssd1 vccd1 vccd1 net1392 _18300__1392/LO sky130_fd_sc_hd__conb_1
X_11411_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[10\] _07326_
+ net2492 vssd1 vssd1 vccd1 vccd1 _07336_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11213__A2 _07096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12391_ net1779 _07798_ _07852_ vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__mux2_1
XANTENNA__12410__A1 _07789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08614__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13040__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11342_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[15\] net509 net359
+ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[11\] vssd1 vssd1 vccd1
+ vccd1 _03398_ sky130_fd_sc_hd__a22o_1
X_14130_ net910 _03992_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[13\]
+ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_30_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__15756__A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11273_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[2\] _07100_ _07129_
+ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[58\] _07233_ vssd1 vssd1
+ vccd1 vccd1 _07234_ sky130_fd_sc_hd__a221o_1
X_14061_ _03911_ _03929_ vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input50_A wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10224_ _05908_ _05992_ net893 vssd1 vssd1 vccd1 vccd1 _06249_ sky130_fd_sc_hd__mux2_1
X_13012_ net270 net2635 net460 vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11495__S net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17820_ clknet_leaf_84_wb_clk_i _03163_ _01516_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08393__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10155_ _04176_ net899 net536 _06179_ _06182_ vssd1 vssd1 vccd1 vccd1 _06183_ sky130_fd_sc_hd__o221a_2
XTAP_TAPCELL_ROW_89_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12611__C _07840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17751_ clknet_leaf_86_wb_clk_i _03094_ _01447_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[61\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold6 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[27\]
+ vssd1 vssd1 vccd1 vccd1 net1420 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12477__A1 _03661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14963_ net1214 vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10086_ net366 _05801_ net517 vssd1 vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16702_ clknet_leaf_163_wb_clk_i _02332_ _00398_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13914_ net1555 net984 _03793_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[28\]
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_85_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17682_ clknet_leaf_91_wb_clk_i _03025_ _01378_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[120\]
+ sky130_fd_sc_hd__dfrtp_1
X_14894_ net1191 vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_50_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16633_ clknet_leaf_10_wb_clk_i _02263_ _00329_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13723__B _06350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13845_ net1471 net579 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[23\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_162_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13215__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16564_ clknet_leaf_127_wb_clk_i _02194_ _00260_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_13776_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[21\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[20\] team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[23\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[22\] vssd1
+ vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__or4_1
XFILLER_0_84_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10988_ _06863_ _06966_ _06967_ net963 vssd1 vssd1 vccd1 vccd1 _06968_ sky130_fd_sc_hd__a211o_1
X_18303_ net1395 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
XFILLER_0_57_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15515_ net1147 vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12727_ _04262_ net563 _03698_ vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__or3_4
X_16495_ clknet_leaf_133_wb_clk_i _02125_ _00191_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14835__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18234_ clknet_leaf_57_wb_clk_i net1467 _01929_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_15446_ net1168 vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12658_ net2958 net341 vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17568__D team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[5\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12401__A1 _07836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11609_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[16\] net994 vssd1
+ vssd1 vccd1 vccd1 _07475_ sky130_fd_sc_hd__and2_2
X_18165_ clknet_leaf_139_wb_clk_i _03468_ _01861_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08605__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15377_ net1192 vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09648__B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12589_ _03610_ net1774 net204 vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17116_ clknet_leaf_158_wb_clk_i _02746_ _00812_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_14328_ net533 _05596_ vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__nor2_1
X_18096_ clknet_leaf_69_wb_clk_i _03419_ _01792_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_29_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwire381 _04342_ vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__buf_4
Xhold406 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[121\] vssd1 vssd1
+ vccd1 vccd1 net1820 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold417 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[72\] vssd1 vssd1
+ vccd1 vccd1 net1831 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10963__A1 _06898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold428 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[14\] vssd1 vssd1
+ vccd1 vccd1 net1842 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold439 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[65\] vssd1 vssd1
+ vccd1 vccd1 net1853 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17047_ clknet_leaf_145_wb_clk_i _02677_ _00743_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14259_ _04035_ _04043_ vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout908 net909 vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__clkbuf_2
Xfanout919 _07367_ vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_74_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[18\]
+ net691 net644 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[18\]
+ _04886_ vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_74_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_146_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1106 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2520 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1117 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net2531 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12468__A1 _07816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1128 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2542 sky130_fd_sc_hd__dlygate4sd3_1
X_08751_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[21\]
+ net816 net788 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[21\]
+ _04821_ vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__a221o_1
X_17949_ clknet_leaf_32_wb_clk_i _03288_ _01645_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1139 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 net2553 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_124_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08682_ _04344_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[23\]
+ _04362_ vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08286__Y _04368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13125__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09097__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09636__A2 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09303_ _04269_ _05307_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_172_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12640__A1 _07816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08844__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12964__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_124_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_63_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1077_A net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09234_ _05284_ vssd1 vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09165_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[11\]
+ net837 net778 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1244_A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08116_ net1028 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[3\]
+ net975 _04207_ vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09096_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[12\]
+ net648 net602 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[12\]
+ _05152_ vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__a221o_1
XFILLER_0_82_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08047_ net1144 vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1032_X net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold940 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2354 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold951 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold973 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2387 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09021__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold984 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net2398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2409 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout492_X net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout871_A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09998_ _06025_ _06026_ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__nand2_1
XANTENNA__12459__A1 _03663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08949_ _04990_ _05011_ vssd1 vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_4_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout757_X net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11960_ _07756_ _07760_ _07757_ vssd1 vssd1 vccd1 vccd1 _07772_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_163_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_174_Left_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10911_ _06219_ _06904_ net956 vssd1 vssd1 vccd1 vccd1 _06905_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout924_X net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11891_ _07665_ _07699_ vssd1 vssd1 vccd1 vccd1 _07703_ sky130_fd_sc_hd__xnor2_2
XANTENNA__09740__C net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13035__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13630_ net1989 net224 net390 vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10842_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[1\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06839_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_80_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12631__A1 _03663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12874__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13561_ net2563 net195 net398 vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10773_ _04166_ team_05_WB.instance_to_wrap.total_design.key_confirm team_05_WB.instance_to_wrap.total_design.key_data
+ vssd1 vssd1 vccd1 vccd1 _06770_ sky130_fd_sc_hd__mux2_1
XANTENNA__08835__B1 _04406_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12727__X _03699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15300_ net1237 vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__inv_2
X_12512_ net1736 _03662_ net209 vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__mux2_1
X_16280_ net1255 vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13492_ net305 net2770 net408 vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15231_ net1180 vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__inv_2
X_12443_ net1732 _03662_ net213 vssd1 vssd1 vccd1 vccd1 _03190_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15162_ net1063 vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__inv_2
X_12374_ net1705 _03657_ net216 vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14113_ _03976_ _03975_ vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__and2b_1
X_11325_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[112\] _07104_
+ _07270_ _07283_ vssd1 vssd1 vccd1 vccd1 _07284_ sky130_fd_sc_hd__a211o_1
XFILLER_0_132_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15093_ net1059 vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_56_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14044_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[10\] _03912_ vssd1
+ vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__xnor2_1
X_11256_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[3\] _07092_ _07129_
+ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[59\] vssd1 vssd1 vccd1
+ vccd1 _07218_ sky130_fd_sc_hd__a22o_1
XANTENNA__13718__B _06445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09012__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17474__Q team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[9\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08366__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10207_ _04554_ net553 _06055_ _05916_ vssd1 vssd1 vccd1 vccd1 _06233_ sky130_fd_sc_hd__o22a_1
XFILLER_0_66_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11187_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[110\] _07102_
+ _07103_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[118\] vssd1
+ vssd1 vccd1 vccd1 _07152_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17803_ clknet_leaf_90_wb_clk_i _03146_ _01499_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[113\]
+ sky130_fd_sc_hd__dfrtp_1
X_10138_ _06164_ _06165_ vssd1 vssd1 vccd1 vccd1 _06166_ sky130_fd_sc_hd__nand2_1
X_15995_ net1128 vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__inv_2
X_17734_ clknet_leaf_87_wb_clk_i _03077_ _01430_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13734__A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10069_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[22\] team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[21\]
+ _06097_ vssd1 vssd1 vccd1 vccd1 _06098_ sky130_fd_sc_hd__and3_1
X_14946_ net1204 vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_141_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17665_ clknet_leaf_98_wb_clk_i _03008_ _01361_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[103\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_141_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14877_ net1089 vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__inv_2
XANTENNA__09650__C net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16616_ clknet_leaf_204_wb_clk_i _02246_ _00312_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13828_ net1509 net578 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[6\]
+ sky130_fd_sc_hd__and2_1
X_17596_ clknet_leaf_51_wb_clk_i _02967_ _01292_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_access
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16547_ clknet_leaf_197_wb_clk_i _02177_ _00243_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13759_ net923 _06907_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[27\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__08826__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12784__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16478_ clknet_leaf_184_wb_clk_i _02108_ _00174_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14284__B _06500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18217_ clknet_leaf_79_wb_clk_i net1524 _01912_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_15429_ net1113 vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18148_ clknet_leaf_176_wb_clk_i _03451_ _01844_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_117_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold203 team_05_WB.instance_to_wrap.total_design.keypad0.key_counter\[3\] vssd1 vssd1
+ vccd1 vccd1 net1617 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_117_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold214 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[34\] vssd1 vssd1
+ vccd1 vccd1 net1628 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18079_ clknet_leaf_85_wb_clk_i _00020_ _01775_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold225 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[101\] vssd1 vssd1
+ vccd1 vccd1 net1639 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold236 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[78\] vssd1 vssd1
+ vccd1 vccd1 net1650 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold247 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[30\] vssd1 vssd1
+ vccd1 vccd1 net1661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[3\] vssd1 vssd1
+ vccd1 vccd1 net1672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[122\] vssd1 vssd1
+ vccd1 vccd1 net1683 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ _05553_ _05949_ _05942_ vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09003__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10149__C1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout705 _04292_ vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__buf_6
XANTENNA__08357__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout716 _04286_ vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__clkbuf_4
Xfanout727 _07355_ vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_165_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09852_ net360 _05879_ vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__nor2_2
Xfanout738 _04421_ vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_165_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout749 net751 vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__clkbuf_8
X_08803_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[19\]
+ net818 net785 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[19\]
+ _04872_ vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__a221o_1
X_09783_ _05809_ _05813_ _05464_ vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__a21bo_1
XANTENNA__12959__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08734_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[21\]
+ net713 net599 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[21\]
+ _04803_ vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_1_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08665_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[23\]
+ net852 net804 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[23\]
+ _04738_ vssd1 vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout452_A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1194_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08596_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[25\]
+ net808 net783 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[25\]
+ _04659_ vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12694__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08817__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout717_A _04286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13810__C net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09217_ _05262_ _05264_ _05266_ _05268_ vssd1 vssd1 vccd1 vccd1 _05269_ sky130_fd_sc_hd__or4_1
XANTENNA__10508__A net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09719__D net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_860 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09148_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[11\]
+ net606 _05191_ net719 vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__a211o_1
XANTENNA__09242__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08596__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09079_ _05131_ _05132_ _05134_ _05136_ vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__or4_1
XFILLER_0_102_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11110_ _07071_ _07073_ _07075_ _07069_ vssd1 vssd1 vccd1 vccd1 _07077_ sky130_fd_sc_hd__a31o_1
XFILLER_0_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_3__f_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_3__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_12090_ _07901_ _07898_ _07893_ vssd1 vssd1 vccd1 vccd1 _07902_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_9_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13877__B1 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold770 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net2184 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout874_X net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold781 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net2195 sky130_fd_sc_hd__dlygate4sd3_1
X_11041_ net1046 _07010_ vssd1 vssd1 vccd1 vccd1 _07011_ sky130_fd_sc_hd__nand2_1
XANTENNA__08348__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold792 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2206 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10155__A2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12869__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14800_ net1093 vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15780_ net1299 vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__inv_2
X_12992_ net321 net2092 net464 vssd1 vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__mux2_1
XANTENNA__09848__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1470 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2884 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1481 net81 vssd1 vssd1 vccd1 vccd1 net2895 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input13_A DAT_I[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14731_ net1070 vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__inv_2
X_11943_ _07730_ _07737_ _07739_ vssd1 vssd1 vccd1 vccd1 _07755_ sky130_fd_sc_hd__and3_1
Xhold1492 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2906 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11655__A2 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17450_ clknet_leaf_46_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[18\]
+ _01146_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08520__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14662_ net1280 vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__inv_2
X_11874_ _07650_ _07672_ _07673_ vssd1 vssd1 vccd1 vccd1 _07686_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_157_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16401_ clknet_leaf_168_wb_clk_i _02031_ _00097_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13613_ net2400 net291 net392 vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__mux2_1
X_17381_ clknet_leaf_60_wb_clk_i net1424 _01077_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10825_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[10\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06822_ sky130_fd_sc_hd__nand2_1
X_14593_ net1219 vssd1 vssd1 vccd1 vccd1 _00223_ sky130_fd_sc_hd__inv_2
X_16332_ net1117 vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13544_ net2686 net276 net403 vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__mux2_1
XANTENNA__09481__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10756_ net362 _05801_ vssd1 vssd1 vccd1 vccd1 _06754_ sky130_fd_sc_hd__or2_1
XANTENNA__17469__Q team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10091__A1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16263_ net1117 vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__inv_2
X_13475_ net259 net2203 net409 vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__mux2_1
X_10687_ _05553_ _05949_ vssd1 vssd1 vccd1 vccd1 _06689_ sky130_fd_sc_hd__xor2_1
X_18002_ clknet_leaf_82_wb_clk_i _03341_ _01698_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15214_ net1187 vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12426_ _03604_ net1827 net215 vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__mux2_1
X_16194_ net1145 vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08587__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13729__A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11040__B1 _06847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12055__D _07478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15145_ net1221 vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12357_ _03648_ _03650_ _03651_ vssd1 vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11308_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[0\] _07100_ _07126_
+ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[80\] vssd1 vssd1 vccd1
+ vccd1 _07267_ sky130_fd_sc_hd__a22o_1
X_15076_ net1205 vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__inv_2
X_12288_ _03578_ _03579_ _03582_ vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__o21a_1
XANTENNA__09645__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14027_ net978 _03895_ _03896_ vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__o21ai_1
X_11239_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[108\] _07111_
+ _07129_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[60\] vssd1 vssd1
+ vccd1 vccd1 _07202_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_71_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12779__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17581__D team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[18\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11536__X _07447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15978_ net1289 vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_160_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09839__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14279__B _06729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17717_ clknet_leaf_91_wb_clk_i _03060_ _01413_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[91\]
+ sky130_fd_sc_hd__dfrtp_1
X_14929_ net1212 vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08511__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08450_ _04522_ _04524_ _04526_ _04528_ vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__or4_1
X_17648_ clknet_leaf_54_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[15\]
+ _01344_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08381_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[30\]
+ net851 net784 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[30\]
+ _04461_ vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__a221o_1
XANTENNA__12367__X _03661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17579_ clknet_leaf_73_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[16\]
+ _01275_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11712__A team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13403__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08293__A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14348__A1 _05078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11431__B team_05_WB.instance_to_wrap.wishbone.curr_state\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09002_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[14\]
+ net696 net650 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09224__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_158_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_158_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08578__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_167_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12543__A _07840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout200_A _06107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout502 net505 vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__clkbuf_2
X_09904_ _04944_ _04966_ vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout513 net515 vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__clkbuf_4
Xfanout524 net525 vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12531__A0 _07798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout546 _07467_ vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09852__A net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input5_A DAT_I[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09835_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[20\]
+ net837 net826 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[20\]
+ _05865_ vssd1 vssd1 vccd1 vccd1 _05866_ sky130_fd_sc_hd__a221o_1
Xfanout557 _04259_ vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__buf_2
Xfanout568 _06774_ vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__clkbuf_4
Xfanout579 net580 vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout667_A _04305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08750__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09571__B net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09766_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[0\]
+ net665 _05796_ net720 vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__a211o_1
X_08717_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[22\]
+ _04366_ net755 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[22\]
+ net855 vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__a221o_1
X_09697_ _05702_ _05720_ _05728_ _05729_ vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__or4_1
XFILLER_0_83_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout834_A net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout455_X net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08502__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08648_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[23\]
+ net701 net645 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout622_X net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08579_ _04648_ _04650_ _04652_ _04654_ vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__or4_1
XANTENNA__12598__A0 _03664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13313__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10610_ _06049_ _06300_ _06308_ _06510_ _06614_ vssd1 vssd1 vccd1 vccd1 _06617_ sky130_fd_sc_hd__o221a_1
XFILLER_0_119_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11590_ team_05_WB.instance_to_wrap.wishbone.curr_state\[1\] net1 vssd1 vssd1 vccd1
+ vccd1 _07471_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10509__Y _06521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14339__A1 _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11270__B1 _07130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10541_ net897 _06551_ vssd1 vssd1 vccd1 vccd1 _06552_ sky130_fd_sc_hd__nor2_1
XANTENNA__14339__B2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[12\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13260_ net324 net2933 net436 vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout991_X net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09215__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10472_ _04158_ _05012_ _06485_ vssd1 vssd1 vccd1 vccd1 _06486_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12211_ _07856_ net500 vssd1 vssd1 vccd1 vccd1 _08023_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_40_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08569__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13191_ net325 net2919 net440 vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__mux2_1
XANTENNA__11573__B2 _07434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12142_ _07953_ vssd1 vssd1 vccd1 vccd1 _07954_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_92_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15764__A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12073_ _07878_ _07882_ _07884_ vssd1 vssd1 vccd1 vccd1 _07885_ sky130_fd_sc_hd__or3_1
X_16950_ clknet_leaf_142_wb_clk_i _02580_ _00646_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1012 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11024_ _06828_ _06829_ _06851_ _06996_ vssd1 vssd1 vccd1 vccd1 _06997_ sky130_fd_sc_hd__a31o_1
X_15901_ net1270 vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__inv_2
X_16881_ clknet_leaf_122_wb_clk_i _02511_ _00577_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12599__S net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15832_ net1272 vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10260__X _06284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15763_ net1302 vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__inv_2
X_12975_ net256 net2573 net464 vssd1 vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14714_ net1056 vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__inv_2
X_17502_ clknet_leaf_109_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[5\]
+ _01198_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11926_ _07734_ _07736_ vssd1 vssd1 vccd1 vccd1 _07738_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15694_ net1159 vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ clknet_leaf_60_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[1\]
+ _01129_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13731__B _05921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14645_ net1059 vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11857_ _07652_ _07662_ _07665_ _07666_ _07667_ vssd1 vssd1 vccd1 vccd1 _07669_ sky130_fd_sc_hd__a32o_1
XFILLER_0_170_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12589__A0 _03610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13223__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15004__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10808_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[17\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[17\]
+ vssd1 vssd1 vccd1 vccd1 _06805_ sky130_fd_sc_hd__and2_1
X_17364_ clknet_leaf_38_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[28\]
+ _01060_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14576_ net1182 vssd1 vssd1 vccd1 vccd1 _00206_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09454__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11788_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[6\] net997 vssd1
+ vssd1 vccd1 vccd1 _07600_ sky130_fd_sc_hd__nand2_2
X_16315_ net1141 vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_136_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11261__B1 _07111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13527_ net2628 net199 net402 vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__mux2_1
X_17295_ clknet_leaf_137_wb_clk_i _02925_ _00991_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10739_ _06470_ net347 vssd1 vssd1 vccd1 vccd1 _06738_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_136_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14843__A net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16246_ net1132 vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__inv_2
X_13458_ net2836 net324 net412 vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17576__D team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12409_ _03651_ net1797 net214 vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16177_ net1158 vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__clkbuf_4
X_13389_ net1985 net329 net421 vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__clkbuf_4
Xoutput127 net127 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__buf_2
XANTENNA__08965__C1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15128_ net1201 vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__inv_2
Xoutput138 net138 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__buf_2
Xoutput149 net149 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15674__A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15059_ net1213 vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__inv_2
XANTENNA__08980__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08717__C1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11707__A team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[11\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08732__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09620_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[2\]
+ net668 net610 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_84 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08288__A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09551_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[3\]
+ net614 net611 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[3\]
+ _05587_ vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__a221o_1
XANTENNA__10330__B _06350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08502_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[27\]
+ net783 net749 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[27\]
+ _04574_ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__a221o_1
X_09482_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[4\]
+ net811 net761 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__a22o_1
XANTENNA__09693__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08433_ _04490_ _04511_ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11442__A net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout248_A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13133__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_747 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08364_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[30\]
+ net649 net630 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[30\]
+ _04435_ vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09445__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08799__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12972__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08295_ net942 net1014 net928 vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout415_A _03727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09566__B net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout203_X net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10345__X _06366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18412__1376 vssd1 vssd1 vccd1 vccd1 _18412__1376/HI net1376 sky130_fd_sc_hd__conb_1
XFILLER_0_103_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout784_A net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08971__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1308 net1309 vssd1 vssd1 vccd1 vccd1 net1308 sky130_fd_sc_hd__buf_4
Xfanout310 net312 vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__clkbuf_2
Xfanout321 net322 vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__clkbuf_2
Xfanout332 _06503_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09582__A team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout343 _07528_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout572_X net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout354 _08023_ vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout951_A _04363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout365 net366 vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13308__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11617__A team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[12\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09818_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[20\]
+ net711 net672 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[20\]
+ _05848_ vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__a221o_1
Xfanout387 _03734_ vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__buf_6
Xfanout398 _03731_ vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_55_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10530__A2 _06540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18322__1414 vssd1 vssd1 vccd1 vccd1 net1414 _18322__1414/LO sky130_fd_sc_hd__conb_1
X_09749_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[0\]
+ net887 net866 net863 vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout837_X net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12760_ _04253_ _04262_ net562 vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__or3_4
XFILLER_0_90_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Left_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11711_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[7\] net997 vssd1
+ vssd1 vccd1 vccd1 _07523_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12691_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[8\] _04251_
+ vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__or2_1
XANTENNA__13043__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14430_ net1062 vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__inv_2
X_11642_ net21 net989 net916 net1624 vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14361_ _04099_ _04133_ _04112_ vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_108_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11573_ net2895 net1005 _07355_ _07434_ vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__a22o_1
XANTENNA__12882__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16100_ net1307 vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__inv_2
Xinput18 DAT_I[24] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13312_ net2551 net270 net428 vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput29 DAT_I[5] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
X_10524_ net897 _06534_ _06535_ _06532_ vssd1 vssd1 vccd1 vccd1 _06536_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_94_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17080_ clknet_leaf_30_wb_clk_i _02710_ _00776_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14292_ _04613_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11498__S net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16031_ net1284 vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__inv_2
XANTENNA__09739__A1 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13243_ net264 net2276 net437 vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10455_ _06308_ _06469_ net371 vssd1 vssd1 vccd1 vccd1 _06470_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_131_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11546__A1 _07422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13174_ net264 net2365 net441 vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10386_ net383 _06404_ vssd1 vssd1 vccd1 vccd1 _06405_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12125_ _07923_ _07927_ _07929_ vssd1 vssd1 vccd1 vccd1 _07937_ sky130_fd_sc_hd__and3_1
XANTENNA__08962__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17982_ clknet_leaf_74_wb_clk_i _03321_ _01678_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__dfrtp_1
XANTENNA__13726__B _06273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12056_ _07525_ _07867_ vssd1 vssd1 vccd1 vccd1 _07868_ sky130_fd_sc_hd__nor2_1
X_16933_ clknet_leaf_181_wb_clk_i _02563_ _00629_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_4_9__f_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11007_ _06822_ _06823_ _06856_ vssd1 vssd1 vccd1 vccd1 _06983_ sky130_fd_sc_hd__a21o_1
XANTENNA__08904__A_N _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16864_ clknet_leaf_129_wb_clk_i _02494_ _00560_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09642__D net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15815_ net1300 vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__inv_2
X_16795_ clknet_leaf_193_wb_clk_i _02425_ _00491_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_172_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15746_ net1288 vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12958_ net310 net2386 net468 vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11909_ _07709_ _07712_ _07720_ _07708_ vssd1 vssd1 vccd1 vccd1 _07721_ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15677_ net1168 vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_138_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12889_ net330 net2658 net477 vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17416_ clknet_leaf_50_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[16\]
+ _01112_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14628_ net1230 vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__inv_2
X_18396_ net913 vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09427__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11234__B1 _07121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17347_ clknet_leaf_40_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[11\]
+ _01043_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_14559_ net1178 vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__inv_2
XANTENNA__12792__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08080_ net1027 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[21\]
+ net969 _04189_ vssd1 vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17278_ clknet_leaf_163_wb_clk_i _02908_ _00974_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10993__C1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14292__B team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[26\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16229_ net1247 vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wire373_X net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08953__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08982_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[15\]
+ net778 net774 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[15\]
+ _05043_ vssd1 vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_143_Right_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11437__A _07349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13128__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09603_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[2\]
+ net877 net862 net857 vssd1 vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_127_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12967__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14748__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_30_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09534_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[3\]
+ _04366_ net837 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[3\]
+ net853 vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__a221o_1
XFILLER_0_167_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09666__B1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09130__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[12\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09465_ net374 _05505_ vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1274_A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08416_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[29\]
+ net818 net751 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09396_ _05426_ _05438_ _05439_ _05440_ vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__or4_2
XFILLER_0_80_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_173_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_173_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_164_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08347_ _04426_ _04427_ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_19_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14483__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout418_X net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_102_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_102_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_62_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08278_ net953 _04360_ _04346_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[21\]
+ sky130_fd_sc_hd__a21o_2
XFILLER_0_22_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10240_ _06003_ _06254_ _06264_ vssd1 vssd1 vccd1 vccd1 _06265_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09197__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout787_X net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08944__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10171_ net524 _06197_ vssd1 vssd1 vccd1 vccd1 _06198_ sky130_fd_sc_hd__nor2_1
XANTENNA__16203__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1105 net1106 vssd1 vssd1 vccd1 vccd1 net1105 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1116 net1119 vssd1 vssd1 vccd1 vccd1 net1116 sky130_fd_sc_hd__buf_4
Xfanout1127 net1177 vssd1 vssd1 vccd1 vccd1 net1127 sky130_fd_sc_hd__buf_2
Xfanout1138 net1139 vssd1 vssd1 vccd1 vccd1 net1138 sky130_fd_sc_hd__buf_4
XANTENNA__09743__C net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1149 net1150 vssd1 vssd1 vccd1 vccd1 net1149 sky130_fd_sc_hd__buf_4
XANTENNA__13038__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13930_ _03801_ _03802_ _03803_ _03804_ vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__and4b_2
XTAP_TAPCELL_ROW_35_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout195 net196 vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13861_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[2\]
+ net560 net576 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[2\]
+ net987 vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_87_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12877__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15600_ net1253 vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12812_ net271 net2824 net484 vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__mux2_1
X_16580_ clknet_leaf_182_wb_clk_i _02210_ _00276_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13792_ net1580 net974 net725 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[3\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_158_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15531_ net1132 vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__inv_2
XANTENNA__09121__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12743_ net268 net2841 net492 vssd1 vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18250_ clknet_leaf_51_wb_clk_i _03479_ _01945_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_15462_ net1160 vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__inv_2
X_12674_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[15\]
+ net339 vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__and2_1
XANTENNA__09409__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ clknet_leaf_122_wb_clk_i _02831_ _00897_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14413_ net1081 vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__inv_2
XANTENNA__11216__B1 _07129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18181_ clknet_leaf_36_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[2\]
+ _01876_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11625_ net1879 net1008 net344 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_12__f_wb_clk_i_X clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15393_ net1235 vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17132_ clknet_leaf_0_wb_clk_i _02762_ _00828_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13501__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14344_ _04096_ _04112_ vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__nor2_1
X_11556_ _07379_ _07465_ vssd1 vssd1 vccd1 vccd1 _07467_ sky130_fd_sc_hd__or2_1
XANTENNA__17477__Q team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[12\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10507_ _05104_ _05963_ vssd1 vssd1 vccd1 vccd1 _06519_ sky130_fd_sc_hd__xor2_1
X_17063_ clknet_leaf_201_wb_clk_i _02693_ _00759_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14275_ net2923 net71 net73 vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_150_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwire585 _05762_ vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__clkbuf_1
X_11487_ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[9\] _07397_ _07345_
+ vssd1 vssd1 vccd1 vccd1 _07398_ sky130_fd_sc_hd__mux2_1
XANTENNA__11021__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16014_ net1112 vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09637__D net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13913__C1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09188__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13226_ _06736_ net351 _03720_ vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_150_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10438_ _06277_ _06355_ _06452_ _06453_ vssd1 vssd1 vccd1 vccd1 _06454_ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08396__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13737__A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08935__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13157_ net323 net1912 net444 vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__mux2_1
X_10369_ _05880_ _05886_ _05976_ vssd1 vssd1 vccd1 vccd1 _06388_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10742__A2 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12108_ _07919_ vssd1 vssd1 vccd1 vccd1 _07920_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17965_ clknet_leaf_108_wb_clk_i _03304_ _01661_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dfrtp_1
X_13088_ net315 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[5\]
+ net455 vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__mux2_1
X_12039_ net919 _07849_ vssd1 vssd1 vccd1 vccd1 _07851_ sky130_fd_sc_hd__nor2_1
X_16916_ clknet_leaf_120_wb_clk_i _02546_ _00612_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13692__A1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17896_ clknet_leaf_104_wb_clk_i _03239_ _01592_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Left_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09360__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16847_ clknet_leaf_138_wb_clk_i _02477_ _00543_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12787__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16778_ clknet_leaf_194_wb_clk_i _02408_ _00474_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_157_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09112__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15729_ net1267 vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_122_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09232__A_N _05256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_0_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_75_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08320__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_114_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_76_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09250_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[9\]
+ net618 net599 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08853__X team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[18\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08201_ _04233_ net958 _04270_ _04154_ _04153_ vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_174_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11207__B1 _07110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10613__A1_N team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09181_ net535 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[11\]
+ sky130_fd_sc_hd__inv_2
X_18379_ net1364 vssd1 vssd1 vccd1 vccd1 la_data_out[27] sky130_fd_sc_hd__buf_2
XFILLER_0_8_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13411__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08132_ _04213_ _04217_ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Left_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_170_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09820__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10430__A1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08063_ net1025 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__and2b_1
XFILLER_0_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18321__1413 vssd1 vssd1 vccd1 vccd1 net1413 _18321__1413/LO sky130_fd_sc_hd__conb_1
XFILLER_0_109_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10770__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08965_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[15\]
+ net660 _05027_ net719 vssd1 vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout482_A net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Left_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08896_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[17\]
+ net774 net763 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_153_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_75_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12697__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14478__A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout747_A _04417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout368_X net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_8__f_wb_clk_i_X clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08476__A _04533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09517_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[10\] _04268_
+ _05555_ vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_91_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout914_A net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11997__A1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[18\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09859__X _05888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09448_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[5\]
+ net848 net762 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05490_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_96_Left_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09379_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[6\]
+ net687 net656 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout702_X net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12726__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13321__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11410_ _07328_ _07335_ vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__nor2_1
X_12390_ net1654 _03604_ _03660_ vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__mux2_1
XANTENNA__09811__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11341_ _04216_ _07286_ net508 vssd1 vssd1 vccd1 vccd1 _07296_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_105_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10246__A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18413__A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14060_ _03927_ _03928_ _03858_ vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__a21o_1
X_11272_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[90\] _07096_
+ _07097_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[34\] _07232_
+ vssd1 vssd1 vccd1 vccd1 _07233_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08378__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13011_ net267 net2932 net460 vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__mux2_1
XANTENNA__08917__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_192_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10223_ net2412 net219 net541 vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_70_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_input43_A wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10154_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[30\] _04238_
+ net895 _06181_ vssd1 vssd1 vccd1 vccd1 _06182_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09590__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12180__B _07690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17750_ clknet_leaf_87_wb_clk_i _03093_ _01446_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[60\]
+ sky130_fd_sc_hd__dfrtp_1
X_14962_ net1238 vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__inv_2
Xhold7 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[6\]
+ vssd1 vssd1 vccd1 vccd1 net1421 sky130_fd_sc_hd__dlygate4sd3_1
X_10085_ _05731_ net366 vssd1 vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__nor2_1
XANTENNA__09342__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16701_ clknet_leaf_110_wb_clk_i _02331_ _00397_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13913_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[28\]
+ net561 net577 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[28\]
+ net988 vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__a221o_1
X_17681_ clknet_leaf_100_wb_clk_i _03024_ _01377_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[119\]
+ sky130_fd_sc_hd__dfrtp_1
X_14893_ net1079 vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_50_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12400__S net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13844_ net1490 net579 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[22\]
+ sky130_fd_sc_hd__and2_1
X_16632_ clknet_leaf_32_wb_clk_i _02262_ _00328_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13426__A1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13775_ _03740_ _03742_ _03745_ _03747_ vssd1 vssd1 vccd1 vccd1 _03748_ sky130_fd_sc_hd__or4_2
X_16563_ clknet_leaf_165_wb_clk_i _02193_ _00259_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10987_ net1045 _06534_ vssd1 vssd1 vccd1 vccd1 _06967_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18302_ net1394 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_100_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15514_ net1149 vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12726_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[7\] _04250_
+ vssd1 vssd1 vccd1 vccd1 _03698_ sky130_fd_sc_hd__or2_1
X_16494_ clknet_leaf_178_wb_clk_i _02124_ _00190_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15445_ net1258 vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__inv_2
X_18233_ clknet_leaf_50_wb_clk_i net1462 _01928_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11811__Y _07623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12657_ team_05_WB.instance_to_wrap.total_design.core.instr_fetch net383 vssd1 vssd1
+ vccd1 vccd1 _03693_ sky130_fd_sc_hd__or2_4
XFILLER_0_154_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13231__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11540__A _07380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11608_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[17\] net994 _07472_
+ net1011 net116 vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__a32o_1
XFILLER_0_4_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15376_ net1195 vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__inv_2
X_18164_ clknet_leaf_173_wb_clk_i _03467_ _01860_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_12588_ _03655_ net1826 net203 vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09648__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17115_ clknet_leaf_190_wb_clk_i _02745_ _00811_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire360 _05860_ vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__buf_4
X_14327_ net374 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[5\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[4\] net373 vssd1
+ vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__a22o_1
X_11539_ _07389_ _07420_ _07446_ vssd1 vssd1 vccd1 vccd1 _07450_ sky130_fd_sc_hd__or3_4
X_18095_ clknet_leaf_68_wb_clk_i _03418_ _01791_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__10156__A _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold407 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[0\] vssd1 vssd1
+ vccd1 vccd1 net1821 sky130_fd_sc_hd__dlygate4sd3_1
Xhold418 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[71\] vssd1 vssd1
+ vccd1 vccd1 net1832 sky130_fd_sc_hd__dlygate4sd3_1
X_17046_ clknet_leaf_150_wb_clk_i _02676_ _00742_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14258_ _04035_ _04038_ _04042_ vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__nor3_2
Xhold429 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[84\] vssd1 vssd1
+ vccd1 vccd1 net1843 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_78_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17584__D team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[21\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08369__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08908__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13209_ net269 net2885 net350 vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__mux2_1
X_14189_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[3\] _07027_
+ vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__or2_1
Xfanout909 _03993_ vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__buf_2
XANTENNA__10715__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[21\]
+ net765 net749 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[21\]
+ _04819_ vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__a221o_1
Xhold1107 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 net2521 sky130_fd_sc_hd__dlygate4sd3_1
X_17948_ clknet_leaf_34_wb_clk_i _03287_ _01644_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[28\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1118 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2532 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1129 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2543 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10479__A1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09333__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08681_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[23\]
+ net592 _04750_ _04754_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[23\]
+ sky130_fd_sc_hd__o22a_4
XANTENNA__10479__B2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17879_ clknet_leaf_76_wb_clk_i _03222_ _01575_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_124_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14298__A net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13406__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08541__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11428__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09302_ _05350_ vssd1 vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_172_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09233_ _05282_ _05283_ vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__nor2_2
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout230_A _06367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout328_A _06705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13141__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09164_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[11\]
+ net814 net802 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08115_ net1027 net2654 vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__and2b_1
XFILLER_0_114_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08072__A2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[25\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09095_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[12\]
+ net683 net621 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__a22o_1
XANTENNA__12980__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1237_A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08046_ team_05_WB.instance_to_wrap.total_design.key_confirm vssd1 vssd1 vccd1 vccd1
+ _04168_ sky130_fd_sc_hd__inv_2
Xclkbuf_4_2__f_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_2__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_102_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold930 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold941 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold952 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2366 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09557__C1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout697_A net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold963 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2377 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13808__C net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold974 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net2388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold996 team_05_WB.instance_to_wrap.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 net2410
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09997_ _05078_ net365 vssd1 vssd1 vccd1 vccd1 _06026_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout864_A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout485_X net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1512_A team_05_WB.instance_to_wrap.CPU_DAT_O\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08780__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08948_ net571 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[16\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[16\] vssd1 vssd1 vccd1
+ vccd1 _05011_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_32_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13656__A1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09324__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13824__B net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08879_ _04357_ _04945_ vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout652_X net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13316__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10910_ net1047 _06245_ _06883_ _06903_ vssd1 vssd1 vccd1 vccd1 _06904_ sky130_fd_sc_hd__a2bb2o_1
X_11890_ _07689_ _07695_ _07697_ _07699_ _07700_ vssd1 vssd1 vccd1 vccd1 _07702_ sky130_fd_sc_hd__a2111o_2
XANTENNA__09740__D net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10841_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[1\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06838_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18408__A net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13560_ net2026 net199 net398 vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__mux2_1
X_10772_ team_05_WB.instance_to_wrap.total_design.core.disable_pc_reg _06768_ vssd1
+ vssd1 vccd1 vccd1 _06769_ sky130_fd_sc_hd__nor2_2
XFILLER_0_66_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12511_ net1622 _03661_ net208 vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13491_ net324 net2769 net408 vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__mux2_1
XANTENNA__13051__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1026 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15230_ net1056 vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__inv_2
X_12442_ net1698 _03661_ net212 vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11198__A2 _07099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15161_ net1057 vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12373_ net1761 _07791_ _07852_ vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__mux2_1
XANTENNA__12890__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14112_ _03975_ _03976_ vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__nand2b_1
X_11324_ _07058_ _07085_ _07084_ _07031_ vssd1 vssd1 vccd1 vccd1 _07283_ sky130_fd_sc_hd__a211o_1
X_15092_ net1074 vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_56_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14043_ net979 _03864_ _03886_ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_56_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11255_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[51\] _07110_
+ _07115_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[59\] _07082_
+ vssd1 vssd1 vccd1 vccd1 _07217_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_128_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1081 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10206_ _06230_ _06231_ net531 vssd1 vssd1 vccd1 vccd1 _06232_ sky130_fd_sc_hd__mux2_1
X_11186_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[30\] _07119_
+ _07121_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[86\] vssd1 vssd1
+ vccd1 vccd1 _07151_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17802_ clknet_leaf_95_wb_clk_i _03145_ _01498_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[112\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08771__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10137_ _04656_ net363 vssd1 vssd1 vccd1 vccd1 _06165_ sky130_fd_sc_hd__nand2_1
X_15994_ net1129 vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__inv_2
XANTENNA__09315__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17733_ clknet_leaf_101_wb_clk_i _03076_ _01429_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13734__B _06729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10068_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[20\] _06096_ vssd1
+ vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__and2_1
XANTENNA__17490__Q team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[25\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14945_ net1228 vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__inv_2
XANTENNA__08523__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17664_ clknet_leaf_93_wb_clk_i _03007_ _01360_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_141_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14876_ net1095 vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__inv_2
XANTENNA__09650__D net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18320__1412 vssd1 vssd1 vccd1 vccd1 net1412 _18320__1412/LO sky130_fd_sc_hd__conb_1
XFILLER_0_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16615_ clknet_leaf_200_wb_clk_i _02245_ _00311_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13827_ net1468 net582 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[5\]
+ sky130_fd_sc_hd__and2_1
X_17595_ clknet_leaf_40_wb_clk_i _02966_ _01291_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.next_next_fetch
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13750__A _05212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13758_ _05212_ _06273_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[26\]
+ sky130_fd_sc_hd__and2_1
X_16546_ clknet_leaf_16_wb_clk_i _02176_ _00242_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17579__D team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[16\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11541__Y _07452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12709_ net272 net2884 net496 vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13689_ net2470 net324 net387 vssd1 vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__mux2_1
X_16477_ clknet_leaf_108_wb_clk_i _02107_ _00173_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14284__C _06521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18216_ clknet_leaf_79_wb_clk_i net1640 _01911_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15428_ net1115 vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11189__A2 _07096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15359_ net1184 vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18147_ clknet_leaf_182_wb_clk_i _03450_ _01843_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10397__B1 _06355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10936__A2 _06320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold204 net125 vssd1 vssd1 vccd1 vccd1 net1618 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold215 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[70\] vssd1 vssd1
+ vccd1 vccd1 net1629 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18078_ clknet_leaf_85_wb_clk_i _00019_ _01774_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold226 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[3\] vssd1 vssd1
+ vccd1 vccd1 net1640 sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[2\] vssd1 vssd1
+ vccd1 vccd1 net1651 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold248 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[66\] vssd1 vssd1
+ vccd1 vccd1 net1662 sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ _05806_ _05948_ _05805_ vssd1 vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__o21ai_2
Xhold259 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[12\] vssd1 vssd1
+ vccd1 vccd1 net1673 sky130_fd_sc_hd__dlygate4sd3_1
X_17029_ clknet_leaf_180_wb_clk_i _02659_ _00725_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout706 _04292_ vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__buf_2
X_09851_ net360 _05879_ vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__nand2b_1
XANTENNA__09554__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout717 _04286_ vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__buf_8
Xfanout728 net730 vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_165_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout739 _04421_ vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__buf_4
XANTENNA__08762__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08802_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[19\]
+ net822 net786 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__a22o_1
X_09782_ _05812_ vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08733_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[21\]
+ net677 net626 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[21\]
+ _04804_ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_1_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08514__B1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13136__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08664_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[23\]
+ net776 net735 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12975__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08595_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[25\]
+ net800 _04670_ net856 vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout445_A net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12828__X _03704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout612_A _04319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09216_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[10\]
+ net790 net782 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[10\]
+ _05267_ vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__a221o_1
XFILLER_0_162_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12377__A1 _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09147_ _05195_ _05197_ _05199_ _05201_ vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout400_X net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09078_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[13\]
+ net837 net764 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[13\]
+ _05135_ vssd1 vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout981_A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08029_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[20\] vssd1
+ vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__inv_2
Xhold760 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 net2174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2185 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold782 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2196 sky130_fd_sc_hd__dlygate4sd3_1
X_11040_ _06834_ _06848_ _06847_ vssd1 vssd1 vccd1 vccd1 _07010_ sky130_fd_sc_hd__a21o_1
XANTENNA__09545__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold793 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net2207 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout867_X net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08753__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13394__X _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12991_ net310 net2307 net464 vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__mux2_1
XANTENNA__09751__C net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1460 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 net2874 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08505__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13046__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11942_ _07730_ _07739_ _07737_ vssd1 vssd1 vccd1 vccd1 _07754_ sky130_fd_sc_hd__a21oi_2
Xhold1471 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 net2885 sky130_fd_sc_hd__dlygate4sd3_1
X_14730_ net1111 vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1482 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2896 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1493 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2907 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_24_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14661_ net1191 vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12885__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11873_ _07672_ _07678_ _07673_ vssd1 vssd1 vccd1 vccd1 _07685_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16400_ clknet_leaf_138_wb_clk_i _02030_ _00096_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13612_ net2291 net278 net392 vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10824_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[11\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06821_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17380_ clknet_leaf_61_wb_clk_i net1447 _01076_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_49_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14592_ net1195 vssd1 vssd1 vccd1 vccd1 _00222_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_862 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16331_ net1116 vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__inv_2
X_13543_ net2120 net272 net400 vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10755_ net2252 net326 net539 vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__mux2_1
XANTENNA__08284__A2 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16262_ net1124 vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13474_ net263 net2525 net408 vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__mux2_1
X_10686_ net2216 net313 net541 vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__mux2_1
XANTENNA__12368__A1 _03661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18001_ clknet_leaf_82_wb_clk_i _03340_ _01697_ vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__dfrtp_1
X_15213_ net1079 vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__inv_2
X_12425_ _03664_ net1817 net214 vssd1 vssd1 vccd1 vccd1 _03205_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16193_ net1145 vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15144_ net1218 vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__inv_2
X_12356_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[28\] net995 _03616_
+ vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__a21o_2
XFILLER_0_106_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13729__B _06185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10705__Y _06706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11307_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[16\] _07125_
+ _07129_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[56\] vssd1 vssd1
+ vccd1 vccd1 _07266_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15075_ net1207 vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__inv_2
X_12287_ _03581_ _03573_ _03574_ vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09645__D net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14026_ net978 _04160_ _03893_ _03894_ vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__o211ai_1
X_11238_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[108\] _07102_
+ _07108_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[92\] _07189_
+ vssd1 vssd1 vccd1 vccd1 _07201_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_71_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12540__A1 _03641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08744__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13745__A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11169_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[47\] _07113_
+ _07118_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[71\] vssd1 vssd1
+ vccd1 vccd1 _07135_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_143_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15977_ net1268 vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_160_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17716_ clknet_leaf_84_wb_clk_i _03059_ _01412_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[90\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14279__C _06743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14928_ net1182 vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17647_ clknet_leaf_70_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[14\]
+ _01343_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14859_ net1075 vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_69_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_920 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08380_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[30\]
+ net754 net749 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17578_ clknet_leaf_73_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[15\]
+ _01274_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16529_ clknet_leaf_172_wb_clk_i _02159_ _00225_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12096__A _07864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08293__B net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09001_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[14\]
+ net702 net604 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08580__Y _04656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08810__A_N net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09903_ net376 _04921_ vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__nand2b_1
Xclkbuf_leaf_198_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_198_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09527__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout503 net505 vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout514 net515 vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout525 _05634_ vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__buf_2
Xfanout536 net538 vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08735__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout395_A _03732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout547 _07466_ vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__buf_4
XFILLER_0_10_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09834_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[20\]
+ net764 net737 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_127_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_127_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10631__X _06637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout558 net561 vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__buf_2
XANTENNA__10542__B1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout569 _06774_ vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__clkbuf_2
X_09765_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[0\]
+ net640 net594 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__a22o_1
XANTENNA__09571__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08716_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[22\]
+ net823 net805 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[22\]
+ _04788_ vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__a221o_1
X_09696_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[1\]
+ net711 _05715_ _05717_ _05719_ vssd1 vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__a2111o_1
X_08647_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[23\]
+ net661 net603 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout350_X net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout827_A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout448_X net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08578_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[25\]
+ net696 net641 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[25\]
+ _04653_ vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10078__X _06107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout615_X net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10540_ _06092_ _06550_ vssd1 vssd1 vccd1 vccd1 _06551_ sky130_fd_sc_hd__or2_1
XANTENNA__14339__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10471_ _05013_ net551 vssd1 vssd1 vccd1 vccd1 _06485_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_157_Right_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12210_ _07856_ net500 vssd1 vssd1 vccd1 vccd1 _08022_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_40_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13190_ net321 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[2\]
+ net440 vssd1 vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__mux2_1
XANTENNA__09766__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09746__C _04287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout984_X net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12141_ _07902_ _07910_ _07952_ vssd1 vssd1 vccd1 vccd1 _07953_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_92_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12072_ net547 _07552_ vssd1 vssd1 vccd1 vccd1 _07884_ sky130_fd_sc_hd__nand2_2
XFILLER_0_25_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold590 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2004 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11325__A2 _07104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15900_ net1302 vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__inv_2
X_11023_ net1045 _06995_ vssd1 vssd1 vccd1 vccd1 _06996_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16880_ clknet_leaf_123_wb_clk_i _02510_ _00576_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_15831_ net1302 vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_32_Left_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15762_ net1297 vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__inv_2
X_12974_ net253 net2881 net464 vssd1 vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__mux2_1
XANTENNA__09151__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1290 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2704 sky130_fd_sc_hd__dlygate4sd3_1
X_17501_ clknet_leaf_114_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[4\]
+ _01197_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_14713_ net1058 vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__inv_2
X_11925_ net549 _07735_ vssd1 vssd1 vccd1 vccd1 _07737_ sky130_fd_sc_hd__nand2_2
X_15693_ net1160 vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__inv_2
XANTENNA_output112_A net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13504__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17432_ clknet_leaf_56_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[0\]
+ _01128_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14644_ net1068 vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__inv_2
X_11856_ _07666_ _07667_ vssd1 vssd1 vccd1 vccd1 _07668_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10807_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[17\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[17\]
+ vssd1 vssd1 vccd1 vccd1 _06804_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17363_ clknet_leaf_34_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[27\]
+ _01059_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14575_ net1233 vssd1 vssd1 vccd1 vccd1 _00205_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08257__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11787_ _07583_ _07586_ _07587_ _07582_ vssd1 vssd1 vccd1 vccd1 _07599_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_64_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16314_ net1124 vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__inv_2
X_10738_ net2653 net321 net539 vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13526_ net557 _03697_ _03707_ vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_136_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08681__X team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[23\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17294_ clknet_leaf_177_wb_clk_i _02924_ _00990_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_41_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16245_ net1124 vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13457_ net2352 net323 net412 vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__mux2_1
X_10669_ _05508_ _05808_ vssd1 vssd1 vccd1 vccd1 _06672_ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12408_ _03662_ net1790 net214 vssd1 vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16176_ net1163 vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__inv_2
X_13388_ net2063 net314 net422 vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__mux2_1
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__clkbuf_4
XANTENNA__12363__B _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__clkbuf_4
XANTENNA__10221__C1 _06243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput128 net128 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__clkbuf_4
X_12339_ _03536_ _03540_ _03517_ _03530_ vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__a211o_1
XFILLER_0_121_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15127_ net1105 vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__inv_2
Xoutput139 net139 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09509__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15058_ net1232 vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12513__A1 _03651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11316__A2 _07099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08717__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14009_ _03852_ _03855_ _03878_ vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__or3b_1
XANTENNA__09672__B net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10524__B1 _06535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08193__A1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09390__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_50_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09017__X _05078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11707__B _07379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08288__B net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09550_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[3\]
+ net704 net632 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_20_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09142__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08501_ _04576_ _04578_ vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_108_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09481_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[4\]
+ net772 net742 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[4\]
+ _05520_ vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__a221o_1
XANTENNA__08496__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13414__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11723__A team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[11\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08432_ net573 _04510_ _04361_ vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11442__B _07354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08363_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[30\]
+ net666 _04443_ net721 vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__a211o_1
XANTENNA__08248__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08294_ _04236_ _04240_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[21\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[20\] _04230_ vssd1
+ vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout408_A _03728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11004__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08956__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08420__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout300 _06621_ vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_111_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout311 net312 vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__buf_2
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1309 net1310 vssd1 vssd1 vccd1 vccd1 net1309 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11307__A2 _07125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12504__A1 _03650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08708__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout398_X net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout322 net323 vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__buf_2
Xfanout333 _06073_ vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10515__B1 _06051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout344 net345 vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__buf_2
Xfanout355 _08023_ vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__buf_1
Xfanout366 net368 vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__buf_2
XANTENNA__09381__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09817_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[20\]
+ net683 net636 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__a22o_1
XANTENNA__10080__Y _06108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout388 _03733_ vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__clkbuf_8
Xfanout399 _03731_ vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__buf_4
X_09748_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[0\]
+ net886 _04287_ net868 vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__and4_1
XANTENNA__08766__X team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[21\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13832__B net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout732_X net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09679_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[1\]
+ net876 net870 net865 vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__and4_1
XANTENNA__08487__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_95_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13324__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1055 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11710_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[8\] net997 vssd1
+ vssd1 vccd1 vccd1 _07522_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12690_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[8\] _04251_
+ vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_24_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11641_ net22 net989 net916 net2926 vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__o22a_1
XFILLER_0_25_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09597__X team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14360_ _04113_ _04131_ _04132_ vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__nand3_1
X_11572_ net1917 net1006 _07355_ _07396_ vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_42_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13311_ net2335 net268 net428 vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__mux2_1
Xinput19 DAT_I[25] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
X_10523_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[14\] net903 net965
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[14\] vssd1 vssd1
+ vccd1 vccd1 _06535_ sky130_fd_sc_hd__a22oi_4
XANTENNA__10451__C1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14291_ _04573_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_94_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13242_ net256 net2360 net436 vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__mux2_1
X_16030_ net1283 vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__inv_2
XANTENNA_input73_A wbs_stb_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09739__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10454_ _06396_ _06468_ net528 vssd1 vssd1 vccd1 vccd1 _06469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13173_ net257 net2049 net441 vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__mux2_1
X_10385_ _06400_ _06403_ vssd1 vssd1 vccd1 vccd1 _06404_ sky130_fd_sc_hd__or2_2
XFILLER_0_58_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10754__B1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_107_Left_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12124_ _07925_ _07934_ _07935_ vssd1 vssd1 vccd1 vccd1 _07936_ sky130_fd_sc_hd__a21bo_1
X_17981_ clknet_leaf_106_wb_clk_i _03320_ _01677_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12055_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[11\] _07379_ _07465_
+ _07478_ vssd1 vssd1 vccd1 vccd1 _07867_ sky130_fd_sc_hd__or4_2
X_16932_ clknet_leaf_183_wb_clk_i _02562_ _00628_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12403__S net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08389__A net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11006_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[11\] net568 _06981_
+ _06982_ vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__a22o_1
X_16863_ clknet_leaf_148_wb_clk_i _02493_ _00559_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_15814_ net1295 vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__inv_2
X_16794_ clknet_leaf_13_wb_clk_i _02424_ _00490_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13742__B _06591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15745_ net1275 vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_29_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12957_ net328 net2739 net469 vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__mux2_1
XANTENNA__08478__A2 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_66_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_116_Left_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13234__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_104_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_59_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11908_ _07710_ _07712_ _07707_ vssd1 vssd1 vccd1 vccd1 _07720_ sky130_fd_sc_hd__a21boi_1
X_15676_ net1168 vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_138_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ net313 net2334 net478 vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17415_ clknet_leaf_60_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[15\]
+ _01111_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10690__C1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14627_ net1203 vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18395_ net913 vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__clkbuf_1
X_11839_ _07625_ _07627_ vssd1 vssd1 vccd1 vccd1 _07651_ sky130_fd_sc_hd__nand2_1
XANTENNA__12431__A0 _03666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10037__A2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17346_ clknet_leaf_42_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[10\]
+ _01042_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14558_ net1056 vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17587__D team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[24\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13509_ net2150 net268 net404 vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17277_ clknet_leaf_128_wb_clk_i _02907_ _00973_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_14489_ net1051 vssd1 vssd1 vccd1 vccd1 _00119_ sky130_fd_sc_hd__inv_2
XANTENNA__08650__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10993__B1 _06898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16228_ net1193 vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08938__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16159_ net1165 vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__inv_2
XANTENNA__08402__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08981_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[15\]
+ net833 net733 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__a22o_1
XANTENNA__11718__A _07379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13409__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08299__A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09363__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire533_X net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_143_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11170__B1 _07119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13933__A _07451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09602_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[2\]
+ net885 net875 net871 vssd1 vssd1 vccd1 vccd1 _05637_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_127_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09115__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09533_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[3\]
+ net786 net778 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[3\]
+ _05562_ vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__a221o_1
XFILLER_0_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08469__A2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout260_A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09666__A1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13144__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09464_ net573 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[5\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[5\] vssd1 vssd1 vccd1
+ vccd1 _05505_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08874__C1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08415_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[29\]
+ net815 net756 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12983__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09395_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[6\]
+ net636 net622 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[6\]
+ _05427_ vssd1 vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout525_A _05634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12422__A0 _03645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09858__A _05886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08346_ net381 _04361_ _04425_ vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08277_ _04152_ _04358_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08641__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout894_A _04279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08929__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15595__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_142_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_142_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_120_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1222_X net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_182_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_131_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10736__B1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10170_ net521 _06195_ _06196_ vssd1 vssd1 vccd1 vccd1 _06197_ sky130_fd_sc_hd__a21o_1
XANTENNA__13827__B net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout682_X net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13319__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1106 net1107 vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__buf_2
Xfanout1117 net1119 vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__buf_4
Xfanout1128 net1130 vssd1 vssd1 vccd1 vccd1 net1128 sky130_fd_sc_hd__buf_4
Xfanout1139 net1141 vssd1 vssd1 vccd1 vccd1 net1139 sky130_fd_sc_hd__buf_4
XANTENNA__09743__D net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout196 _06184_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__buf_1
X_13860_ net1513 net982 _03766_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[1\]
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_87_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09106__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13989__B1 _07451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12811_ net267 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[16\]
+ net484 vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__mux2_1
X_13791_ net1716 net972 net726 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[2\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_96_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_754 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13054__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15530_ net1149 vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__inv_2
X_12742_ net259 net2503 net493 vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10672__C1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15461_ net1171 vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12673_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[16\]
+ net339 vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__and2_1
XANTENNA__12893__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17200_ clknet_leaf_124_wb_clk_i _02830_ _00896_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14412_ net1109 vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__inv_2
X_11624_ net2642 net1008 net344 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__a22o_1
X_18180_ clknet_leaf_38_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[1\]
+ _01875_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15392_ net1197 vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_133_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17131_ clknet_leaf_188_wb_clk_i _02761_ _00827_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11555_ _07379_ _07465_ vssd1 vssd1 vccd1 vccd1 _07466_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14343_ _04097_ _04098_ _04113_ _04114_ vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__and4_1
XFILLER_0_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08632__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10506_ net2702 net271 net539 vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__mux2_1
X_14274_ net985 net574 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.next_read
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_150_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17062_ clknet_leaf_117_wb_clk_i _02692_ _00758_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11486_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[9\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[9\]
+ net1034 vssd1 vssd1 vccd1 vccd1 _07397_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_150_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire586 _05759_ vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__buf_1
XANTENNA__13913__B1 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16013_ net1112 vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__inv_2
X_13225_ net2951 net351 vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__nand2_1
X_10437_ _04925_ _06056_ vssd1 vssd1 vccd1 vccd1 _06453_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13156_ net309 net2902 net444 vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__mux2_1
X_10368_ _05886_ _06386_ vssd1 vssd1 vccd1 vccd1 _06387_ sky130_fd_sc_hd__xnor2_4
X_12107_ _07915_ _07916_ _07918_ vssd1 vssd1 vccd1 vccd1 _07919_ sky130_fd_sc_hd__a21o_1
XANTENNA__11538__A _07379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13087_ net317 net2667 net452 vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__mux2_1
X_17964_ clknet_leaf_107_wb_clk_i _03303_ _01660_ vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__dfrtp_1
X_10299_ net893 _06320_ vssd1 vssd1 vccd1 vccd1 _06321_ sky130_fd_sc_hd__or2_1
X_12038_ _07847_ _07849_ _07844_ vssd1 vssd1 vccd1 vccd1 _07850_ sky130_fd_sc_hd__a21o_1
X_16915_ clknet_leaf_167_wb_clk_i _02545_ _00611_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_17895_ clknet_leaf_89_wb_clk_i _03238_ _01591_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08699__A2 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13753__A net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16846_ clknet_leaf_170_wb_clk_i _02476_ _00542_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16777_ clknet_leaf_21_wb_clk_i _02407_ _00473_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13989_ team_05_WB.instance_to_wrap.CPU_DAT_O\[5\] net546 _07451_ vssd1 vssd1 vccd1
+ vccd1 _03860_ sky130_fd_sc_hd__a21o_1
XFILLER_0_149_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15728_ net1272 vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_157_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09949__Y _05978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15659_ net1248 vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_174_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08871__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08200_ _04233_ net958 _04270_ _04156_ _04155_ vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_174_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09180_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[11\]
+ net590 _05227_ _05233_ vssd1 vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__o22ai_4
XTAP_TAPCELL_ROW_174_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18378_ net1363 vssd1 vssd1 vccd1 vccd1 la_data_out[26] sky130_fd_sc_hd__buf_2
XFILLER_0_44_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08131_ _04213_ _04217_ vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__nor2_1
XFILLER_0_133_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17329_ clknet_leaf_118_wb_clk_i _02959_ _01025_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_170_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08623__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08062_ net1024 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[30\]
+ net969 _04180_ vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__a22o_1
XANTENNA__10430__A2 _06445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_1__f_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_1__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10718__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13380__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13139__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08964_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[15\]
+ net621 net617 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05027_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1015_A _04347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09336__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12978__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08895_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[17\]
+ net840 net759 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout475_A _03706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12891__A0 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout642_A net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12643__A0 _03641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09516_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[15\] net966
+ _04267_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[23\] _05554_
+ vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09447_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[5\]
+ net784 net780 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[5\]
+ _05488_ vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout430_X net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08862__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13602__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09378_ _05420_ _05421_ vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__or2_2
XFILLER_0_47_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08329_ net1015 net948 net928 vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__and3_1
XFILLER_0_151_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08614__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11340_ _07287_ _07291_ _07294_ vssd1 vssd1 vccd1 vccd1 _07295_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_132_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10246__B _06270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout897_X net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11271_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[114\] _07103_
+ _07124_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[26\] _07231_
+ vssd1 vssd1 vccd1 vccd1 _07232_ sky130_fd_sc_hd__a221o_1
XFILLER_0_15_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13010_ net259 net2905 net461 vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__mux2_1
X_10222_ net383 _06247_ vssd1 vssd1 vccd1 vccd1 _06248_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_37_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13049__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10153_ _06103_ _06180_ vssd1 vssd1 vccd1 vccd1 _06181_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_101_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_89_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09327__B1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input36_A gpio_in[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14961_ net1216 vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_54_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10084_ net523 net366 vssd1 vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__and2_1
XANTENNA__12888__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1422 sky130_fd_sc_hd__dlygate4sd3_1
X_16700_ clknet_leaf_161_wb_clk_i _02330_ _00396_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13912_ net1537 net983 _03792_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[27\]
+ sky130_fd_sc_hd__o21a_1
X_17680_ clknet_leaf_104_wb_clk_i _03023_ _01376_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[118\]
+ sky130_fd_sc_hd__dfrtp_1
X_14892_ net1071 vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__inv_2
X_16631_ clknet_leaf_146_wb_clk_i _02261_ _00327_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13843_ net1485 net579 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[21\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_18_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16562_ clknet_leaf_127_wb_clk_i _02192_ _00258_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13774_ _03743_ _03744_ _03746_ vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__or3_1
X_10986_ _06812_ _06862_ net1045 vssd1 vssd1 vccd1 vccd1 _06966_ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18301_ net1393 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
XFILLER_0_57_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15513_ net1161 vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12725_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[7\] _04250_
+ vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__nor2_1
X_16493_ clknet_leaf_160_wb_clk_i _02123_ _00189_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08853__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13512__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18232_ clknet_leaf_50_wb_clk_i net1478 _01927_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_15444_ net1258 vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_152_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12656_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[11\] _04249_
+ team_05_WB.instance_to_wrap.total_design.core.instr_fetch vssd1 vssd1 vccd1 vccd1
+ _03692_ sky130_fd_sc_hd__a21o_1
XFILLER_0_167_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11607_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[18\] net994 _07472_
+ net1011 net117 vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__a32o_1
X_18163_ clknet_leaf_114_wb_clk_i _03466_ _01859_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_12587_ _03646_ net1927 _03681_ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15375_ net1283 vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__inv_2
XANTENNA__08605__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09648__D net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17114_ clknet_leaf_12_wb_clk_i _02744_ _00810_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_14326_ net535 _05208_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[12\]
+ _05165_ vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__o2bb2a_1
X_18094_ clknet_leaf_68_wb_clk_i _03417_ _01790_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_11538_ _07379_ _07447_ vssd1 vssd1 vccd1 vccd1 _07449_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10156__B _06183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold408 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[53\] vssd1 vssd1
+ vccd1 vccd1 net1822 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13748__A net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold419 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[43\] vssd1 vssd1
+ vccd1 vccd1 net1833 sky130_fd_sc_hd__dlygate4sd3_1
X_17045_ clknet_leaf_21_wb_clk_i _02675_ _00741_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_14257_ _00030_ _00029_ _04041_ vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__or3_1
X_11469_ _07369_ _07378_ vssd1 vssd1 vccd1 vccd1 _07380_ sky130_fd_sc_hd__or2_4
XFILLER_0_150_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13208_ _06479_ net2295 net351 vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__mux2_1
X_14188_ _07027_ net729 _03996_ vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__and3b_1
XFILLER_0_1_979 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09030__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13139_ net253 net2875 net444 vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__mux2_1
XANTENNA__10596__A2_N net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14311__B1 _04818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17947_ clknet_leaf_34_wb_clk_i _03286_ _01643_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1108 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2522 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1119 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 net2533 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12798__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08680_ _04739_ _04741_ _04752_ _04753_ vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__or4_1
XFILLER_0_174_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17878_ clknet_leaf_76_wb_clk_i _03221_ _01574_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_124_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14298__B team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[24\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16829_ clknet_leaf_131_wb_clk_i _02459_ _00525_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08829__C1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09097__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09301_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[8\]
+ net718 _05346_ _05349_ vssd1 vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__o22a_4
XFILLER_0_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12386__X _03663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08844__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09232_ _05256_ _05280_ vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__and2b_1
XANTENNA__13422__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09163_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[11\]
+ net822 net806 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__a22o_1
X_08114_ net1032 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[4\]
+ net976 _04206_ vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09094_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[12\]
+ net625 net606 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[12\]
+ _05148_ vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__a221o_1
XANTENNA__11600__B2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[24\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08045_ team_05_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold920 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold931 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold942 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2356 sky130_fd_sc_hd__dlygate4sd3_1
Xhold953 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2367 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold964 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 net2378 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09021__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09574__C net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold975 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 net2389 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout592_A _04368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold986 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2400 sky130_fd_sc_hd__dlygate4sd3_1
Xhold997 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 net2411 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10082__A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09996_ _05034_ net364 vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout1018_X net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09309__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08947_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[16\]
+ net590 _05006_ _05010_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[16\]
+ sky130_fd_sc_hd__o22a_4
XTAP_TAPCELL_ROW_32_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout857_A net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout478_X net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12501__S net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08878_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[17\] _04356_
+ vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_4_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout645_X net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12616__A0 _03651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10840_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[2\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06837_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_80_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10771_ net1042 net961 vssd1 vssd1 vccd1 vccd1 _06768_ sky130_fd_sc_hd__nor2_4
XFILLER_0_17_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08296__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout812_X net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08835__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13332__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12510_ net1975 net500 _03676_ vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13490_ net322 net2807 net408 vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__mux2_1
XANTENNA__09749__C net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12441_ net1616 net500 net212 vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12372_ net1608 _07789_ _07852_ vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__mux2_1
X_15160_ net1244 vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__inv_2
X_11323_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[56\] _07115_
+ _07116_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[72\] _07271_
+ vssd1 vssd1 vccd1 vccd1 _07282_ sky130_fd_sc_hd__a221o_1
X_14111_ _03955_ _03965_ _03968_ vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_132_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15091_ net1217 vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09548__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11254_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[43\] _07113_
+ _07116_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[75\] _07215_
+ vssd1 vssd1 vccd1 vccd1 _07216_ sky130_fd_sc_hd__a221o_1
X_14042_ team_05_WB.instance_to_wrap.CPU_DAT_O\[7\] net546 _07451_ vssd1 vssd1 vccd1
+ vccd1 _03911_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_56_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09012__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10205_ _06166_ _06175_ net520 vssd1 vssd1 vccd1 vccd1 _06231_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11185_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[62\] _07115_
+ _07118_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[70\] vssd1 vssd1
+ vccd1 vccd1 _07150_ sky130_fd_sc_hd__a22o_1
X_17801_ clknet_leaf_100_wb_clk_i _03144_ _01497_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[111\]
+ sky130_fd_sc_hd__dfrtp_1
X_10136_ _04613_ net368 vssd1 vssd1 vccd1 vccd1 _06164_ sky130_fd_sc_hd__nand2_1
X_15993_ net1128 vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_145_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13507__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17732_ clknet_leaf_93_wb_clk_i _03075_ _01428_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12411__S _03667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10067_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[19\] team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[18\]
+ _06095_ vssd1 vssd1 vccd1 vccd1 _06096_ sky130_fd_sc_hd__and3_1
X_14944_ net1102 vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17663_ clknet_leaf_88_wb_clk_i _03006_ _01359_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[101\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_141_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14875_ net1176 vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_141_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11027__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload1_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12607__A0 _03650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16614_ clknet_leaf_119_wb_clk_i _02244_ _00310_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13826_ net1497 net581 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[4\]
+ sky130_fd_sc_hd__and2_1
X_17594_ clknet_leaf_109_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[31\]
+ _01290_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13750__B _06445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16545_ clknet_leaf_151_wb_clk_i _02175_ _00241_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13757_ net923 _06918_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[25\]
+ sky130_fd_sc_hd__nor2_1
X_10969_ _06952_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[18\] net564
+ vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__mux2_1
XANTENNA__10719__X _06720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08826__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13242__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12708_ net268 net2730 net496 vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__mux2_1
X_16476_ clknet_leaf_161_wb_clk_i _02106_ _00172_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13688_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[2\]
+ net322 net387 vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__mux2_1
X_18215_ clknet_leaf_78_wb_clk_i net1978 _01910_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15427_ net1114 vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12639_ net1643 _07821_ _03682_ vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11043__C1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18146_ clknet_leaf_198_wb_clk_i _03449_ _01842_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_15358_ net1065 vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__inv_2
XANTENNA__10397__A1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09251__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11594__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold205 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[19\] vssd1 vssd1
+ vccd1 vccd1 net1619 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_117_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14309_ _04070_ _04078_ _04081_ _04069_ vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__or4b_2
X_18077_ clknet_leaf_84_wb_clk_i _00018_ _01773_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09675__B net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold216 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[99\] vssd1 vssd1
+ vccd1 vccd1 net1630 sky130_fd_sc_hd__dlygate4sd3_1
X_15289_ net1057 vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__inv_2
Xhold227 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[73\] vssd1 vssd1
+ vccd1 vccd1 net1641 sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[22\] vssd1 vssd1
+ vccd1 vccd1 net1652 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09539__B1 _05556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold249 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[102\] vssd1 vssd1
+ vccd1 vccd1 net1663 sky130_fd_sc_hd__dlygate4sd3_1
X_17028_ clknet_leaf_181_wb_clk_i _02658_ _00724_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09003__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09850_ net571 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[20\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[20\] vssd1 vssd1 vccd1
+ vccd1 _05879_ sky130_fd_sc_hd__a21oi_1
Xfanout707 net710 vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__buf_6
XFILLER_0_42_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout718 _04286_ vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__clkbuf_8
Xfanout729 net730 vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_165_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[19\]
+ net845 net778 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[19\]
+ _04870_ vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__a221o_1
X_09781_ _05464_ _05811_ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11726__A _07379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13417__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08732_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[21\]
+ net705 net680 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08663_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[23\]
+ net828 net758 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08594_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[25\]
+ net750 net747 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_138_Right_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08817__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout340_A _03693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1082_A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13152__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout438_A _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10624__A2 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09569__C net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09215_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[10\]
+ net810 net760 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__a22o_1
XANTENNA__12991__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout605_A _04321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09866__A net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09146_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[11\]
+ net652 net614 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[11\]
+ _05200_ vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09242__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09077_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[13\]
+ net844 net768 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__a22o_1
XANTENNA__09585__B net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_49_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08028_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[21\] vssd1
+ vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__inv_2
Xhold750 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2164 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout974_A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold761 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 net2175 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout595_X net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold772 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net2186 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold783 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2197 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold794 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net2208 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10560__A1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[12\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout762_X net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09979_ _06006_ _06007_ vssd1 vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__nand2_1
XANTENNA__13327__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12990_ net328 net2601 net466 vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09751__D net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1450 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2864 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1461 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 net2875 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11941_ _07752_ vssd1 vssd1 vccd1 vccd1 _07753_ sky130_fd_sc_hd__inv_2
Xhold1472 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2886 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1483 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 net2897 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1494 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2908 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14660_ net1229 vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__inv_2
X_11872_ _07597_ _07683_ _07529_ vssd1 vssd1 vccd1 vccd1 _07684_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13611_ net2022 net282 net393 vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__mux2_1
X_10823_ _06819_ vssd1 vssd1 vccd1 vccd1 _06820_ sky130_fd_sc_hd__inv_2
XANTENNA__12065__A1 _07478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10686__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08808__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14591_ net1178 vssd1 vssd1 vccd1 vccd1 _00221_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13062__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16330_ net1118 vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__inv_2
X_13542_ net2175 net269 net400 vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__mux2_1
X_10754_ _06751_ _06752_ net383 vssd1 vssd1 vccd1 vccd1 _06753_ sky130_fd_sc_hd__o21a_1
XANTENNA__09481__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13014__A0 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16261_ net1123 vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_45_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13473_ net257 net2251 net409 vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__mux2_1
X_10685_ _04264_ _06687_ vssd1 vssd1 vccd1 vccd1 _06688_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18000_ clknet_leaf_63_wb_clk_i _03339_ _01696_ vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11025__C1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15212_ net1071 vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__inv_2
XFILLER_0_164_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12424_ net1668 _03663_ _03667_ vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16192_ net1145 vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_97_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15143_ net1199 vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__inv_2
XANTENNA__12406__S net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12355_ _03511_ _03524_ _03528_ _03649_ vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__a31o_2
XFILLER_0_51_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08441__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11306_ net1887 net732 _07265_ vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__o21a_1
X_12286_ _03568_ _03573_ vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__nand2b_1
X_15074_ net1226 vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_147_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11237_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[60\] _07115_
+ _07117_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[52\] _07199_
+ vssd1 vssd1 vccd1 vccd1 _07200_ sky130_fd_sc_hd__a221o_1
X_14025_ _03893_ _03894_ _04160_ vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_112_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13745__B _06540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11168_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[111\] _07102_
+ _07126_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[87\] _07131_
+ vssd1 vssd1 vccd1 vccd1 _07134_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_143_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13237__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10119_ _06145_ _06146_ vssd1 vssd1 vccd1 vccd1 _06147_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_93_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11099_ _04162_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[3\]
+ _07054_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[5\] vssd1
+ vssd1 vccd1 vccd1 _07066_ sky130_fd_sc_hd__o31a_1
X_15976_ net1265 vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__inv_2
XANTENNA__10450__A net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17715_ clknet_leaf_80_wb_clk_i _03058_ _01411_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[89\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_160_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14279__D _06756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14927_ net1280 vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__inv_2
XANTENNA__14857__A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18379__1364 vssd1 vssd1 vccd1 vccd1 _18379__1364/HI net1364 sky130_fd_sc_hd__conb_1
XANTENNA__13761__A net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17646_ clknet_leaf_70_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[13\]
+ _01342_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_14858_ net1122 vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__inv_2
XANTENNA__08855__A net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13809_ net1558 net970 net723 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[20\]
+ sky130_fd_sc_hd__and3_1
X_17577_ clknet_leaf_113_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[14\]
+ _01273_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14789_ net1191 vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__inv_2
XANTENNA__10449__X _06464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16528_ clknet_leaf_167_wb_clk_i _02158_ _00224_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08293__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16459_ clknet_leaf_188_wb_clk_i _02089_ _00155_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_09000_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[14\]
+ net713 net638 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[14\]
+ _05060_ vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__a221o_1
XANTENNA__13556__A1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09224__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11567__B1 _07354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18129_ clknet_leaf_48_wb_clk_i _00025_ _01825_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_167_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09902_ _04880_ _04881_ vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__nor2_2
XFILLER_0_1_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout504 net505 vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout515 _05700_ vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_158_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout526 net527 vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__clkbuf_4
Xfanout537 net538 vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__clkbuf_4
X_09833_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[20\]
+ net802 net774 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[20\]
+ _05862_ vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__a221o_1
Xfanout548 _07449_ vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__buf_2
Xfanout559 net560 vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__buf_2
XANTENNA__10542__A1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10542__B2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13147__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_A _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1026 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09764_ _05791_ _05792_ _05793_ _05794_ vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__or4_1
XANTENNA__09571__D net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_167_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_167_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08715_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[22\]
+ net831 net815 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__a22o_1
XANTENNA__08499__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12986__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09695_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[1\]
+ net672 _05705_ _05709_ _05713_ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_69_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout555_A net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14767__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_99_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08646_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[23\]
+ net693 net674 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08577_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[25\]
+ net708 net673 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout722_A _04285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13821__D _03748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09463__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout510_X net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11270__A2 _07123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08671__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1252_X net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout608_X net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13610__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10470_ net892 _06481_ _06483_ vssd1 vssd1 vccd1 vccd1 _06484_ sky130_fd_sc_hd__o21a_1
XFILLER_0_134_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09215__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09129_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[12\]
+ net590 _05180_ _05184_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[12\]
+ sky130_fd_sc_hd__o22a_4
XFILLER_0_44_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09746__D net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08974__A1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[27\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12140_ _07903_ _07951_ vssd1 vssd1 vccd1 vccd1 _07952_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_1091 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout977_X net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12071_ _07878_ _07882_ vssd1 vssd1 vccd1 vccd1 _07883_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold580 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net1994 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold591 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 net2005 sky130_fd_sc_hd__dlygate4sd3_1
X_11022_ _06828_ _06829_ _06851_ vssd1 vssd1 vccd1 vccd1 _06995_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13057__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15830_ net1263 vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15761_ net1276 vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__inv_2
X_12973_ net247 net2699 net466 vssd1 vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__mux2_1
XANTENNA__12896__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1280 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net2694 sky130_fd_sc_hd__dlygate4sd3_1
X_17500_ clknet_leaf_113_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[3\]
+ _01196_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[3\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold1291 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2705 sky130_fd_sc_hd__dlygate4sd3_1
X_14712_ net1244 vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__inv_2
X_11924_ net549 _07735_ vssd1 vssd1 vccd1 vccd1 _07736_ sky130_fd_sc_hd__and2_1
X_15692_ net1169 vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17431_ clknet_leaf_57_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[31\]
+ _01127_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14643_ net1215 vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11813__B _07623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10269__X _06293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11855_ _07619_ _07628_ _07632_ vssd1 vssd1 vccd1 vccd1 _07667_ sky130_fd_sc_hd__nand3_1
X_10806_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[18\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06803_ sky130_fd_sc_hd__or2_1
X_17362_ clknet_leaf_36_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[26\]
+ _01058_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_99_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14574_ net1187 vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09454__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11786_ _07583_ _07586_ _07587_ _07589_ vssd1 vssd1 vccd1 vccd1 _07598_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_64_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16313_ net1124 vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13525_ net2568 net307 net407 vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__mux2_1
XANTENNA__11261__A2 _07109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17293_ clknet_leaf_162_wb_clk_i _02923_ _00989_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10737_ _04264_ _06736_ vssd1 vssd1 vccd1 vccd1 _06737_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_136_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13520__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16244_ net1131 vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__inv_2
X_13456_ net1990 net311 net413 vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__mux2_1
XANTENNA__17496__Q team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[31\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10668_ net2482 net319 net540 vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12407_ _03661_ net1795 net215 vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16175_ net1153 vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_114_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08414__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13387_ net1973 net318 net421 vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__mux2_1
X_10599_ net2157 net289 net539 vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__mux2_1
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15126_ net1085 vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__inv_2
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__buf_2
X_12338_ _03531_ _03540_ _03536_ vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__a21o_1
Xoutput129 net129 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13756__A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15057_ net1192 vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__inv_2
X_12269_ _07968_ _07977_ _03558_ _03561_ _03562_ vssd1 vssd1 vccd1 vccd1 _03564_ sky130_fd_sc_hd__a32o_1
X_14008_ _03852_ _03855_ _03878_ vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_162_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10524__A1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_133_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09672__C net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08202__X _04285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11707__C _07447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08288__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15959_ net1302 vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__inv_2
X_08500_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[27\]
+ net834 net739 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[27\]
+ _04577_ vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__a221o_1
X_09480_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[4\]
+ net830 net769 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__a22o_1
XANTENNA__09693__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08431_ _04510_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[29\]
+ sky130_fd_sc_hd__inv_2
X_17629_ clknet_leaf_51_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.next_state\[0\]
+ _01325_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.state\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_08362_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[30\]
+ net642 net595 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09445__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09903__A_N net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08653__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08293_ net948 net938 net931 vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13430__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10460__B1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08405__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_172_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1045_A net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09566__D net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16042__A net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1212_A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout301 _06621_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__buf_1
Xfanout312 _06720_ vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__clkbuf_2
Xfanout323 _06737_ vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__buf_2
Xfanout334 _06073_ vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__buf_2
XANTENNA__10515__A1 _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout672_A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09582__C net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout345 net346 vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__buf_2
Xfanout356 _07516_ vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__buf_2
X_09816_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[20\]
+ net656 net632 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[20\]
+ _05846_ vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__a221o_1
Xfanout367 net368 vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__buf_2
XANTENNA__10090__A _05442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout389 _03733_ vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__buf_4
X_09747_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[0\]
+ net886 net875 net861 vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout460_X net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13605__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09678_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[1\]
+ net876 net869 net857 vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__and4_1
X_08629_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[24\]
+ net830 net739 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08892__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout725_X net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11640_ net23 net989 net916 net2857 vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__o22a_1
XFILLER_0_64_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11571_ net1902 net1004 net727 _07407_ vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_42_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08644__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13340__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_64_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13310_ net2348 net261 net431 vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__mux2_1
X_10522_ _06093_ _06533_ vssd1 vssd1 vccd1 vccd1 _06534_ sky130_fd_sc_hd__or2_2
X_14290_ net899 net921 _05921_ _04063_ _06772_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.next_instr_wait
+ sky130_fd_sc_hd__a221oi_1
XFILLER_0_123_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09757__C net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13241_ net253 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[20\]
+ net436 vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__mux2_1
X_10453_ _06429_ _06467_ net518 vssd1 vssd1 vccd1 vccd1 _06468_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_131_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18378__1363 vssd1 vssd1 vccd1 vccd1 _18378__1363/HI net1363 sky130_fd_sc_hd__conb_1
XANTENNA_input66_A wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10384_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[21\] net903 net967
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[21\] _06402_ vssd1
+ vssd1 vccd1 vccd1 _06403_ sky130_fd_sc_hd__a221o_1
X_13172_ net253 net2815 net440 vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12123_ _07923_ _07925_ _07929_ vssd1 vssd1 vccd1 vccd1 _07935_ sky130_fd_sc_hd__or3_1
X_17980_ clknet_leaf_74_wb_clk_i _03319_ _01676_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12054_ _07865_ vssd1 vssd1 vccd1 vccd1 _07866_ sky130_fd_sc_hd__inv_2
X_16931_ clknet_leaf_198_wb_clk_i _02561_ _00627_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11005_ net963 _06572_ net568 vssd1 vssd1 vccd1 vccd1 _06982_ sky130_fd_sc_hd__a21oi_1
X_16862_ clknet_leaf_162_wb_clk_i _02492_ _00558_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_15813_ net1290 vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__inv_2
Xfanout890 net891 vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__buf_2
X_16793_ clknet_leaf_15_wb_clk_i _02423_ _00489_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13515__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15744_ net1264 vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__inv_2
X_12956_ net314 net2240 net470 vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11907_ _07684_ _07714_ _07717_ _07718_ vssd1 vssd1 vccd1 vccd1 _07719_ sky130_fd_sc_hd__or4_1
XFILLER_0_158_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15675_ net1166 vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ net317 net2669 net477 vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__mux2_1
XANTENNA__08883__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17414_ clknet_leaf_60_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[14\]
+ _01110_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_138_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14626_ net1204 vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18394_ net915 vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__clkbuf_1
X_11838_ _07649_ _07644_ _07645_ vssd1 vssd1 vccd1 vccd1 _07650_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09427__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10159__B _06185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17345_ clknet_4_5__leaf_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[9\]
+ _01041_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11234__A2 _07118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ net1090 vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__inv_2
XANTENNA__08635__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11769_ _07567_ _07571_ _07563_ _07564_ vssd1 vssd1 vccd1 vccd1 _07581_ sky130_fd_sc_hd__o211ai_1
XANTENNA__13250__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13508_ net2418 net260 net404 vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__mux2_1
X_17276_ clknet_leaf_157_wb_clk_i _02906_ _00972_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14488_ net1244 vssd1 vssd1 vccd1 vccd1 _00118_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_0__f_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_0__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_16227_ net1227 vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__inv_2
XANTENNA__15966__A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13439_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[20\]
+ net252 net412 vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16158_ net1175 vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09060__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17954__Q net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15109_ net1194 vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__inv_2
X_16089_ net1308 vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__inv_2
X_08980_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[15\]
+ net786 net764 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[15\]
+ _05037_ vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__a221o_1
XANTENNA__10903__A _04170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12498__A1 _07797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11718__B _07447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08299__B net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09601_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[2\]
+ net886 net863 net859 vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__and4_1
XFILLER_0_39_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13425__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09532_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[3\]
+ net844 net818 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[3\]
+ _05561_ vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09666__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09463_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[5\]
+ net593 _05500_ _05504_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[5\]
+ sky130_fd_sc_hd__o22a_4
XFILLER_0_93_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10681__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09698__X _05731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08414_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[29\]
+ net846 net761 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[29\]
+ _04493_ vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09394_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[6\]
+ net695 net633 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[6\]
+ _05429_ vssd1 vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11225__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08626__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08345_ _04361_ _04425_ net381 vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout420_A net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1162_A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout518_A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08276_ _04358_ vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09577__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10085__A _05731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14780__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09874__A _04656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09051__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10736__B2 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout887_A _04281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12504__S net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12489__A1 _03614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_182_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_182_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout1107 net1108 vssd1 vssd1 vccd1 vccd1 net1107 sky130_fd_sc_hd__clkbuf_4
Xfanout1118 net1119 vssd1 vssd1 vccd1 vccd1 net1118 sky130_fd_sc_hd__buf_2
Xfanout1129 net1130 vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout675_X net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_111_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_111_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_156_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout197 net200 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout842_X net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13335__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12810_ net261 net2370 net485 vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__mux2_1
X_13790_ net1562 net975 net726 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[1\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__09657__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ net263 net2292 net492 vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08865__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14955__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15460_ net1167 vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__inv_2
X_12672_ net2613 net340 vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__and2_1
XFILLER_0_132_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09409__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ net1070 vssd1 vssd1 vccd1 vccd1 _00041_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ net1930 net1009 net344 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__a22o_1
XANTENNA__12413__A1 _07793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11216__A2 _07108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15391_ net1182 vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__inv_2
XANTENNA__08617__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13070__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10424__B1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17130_ clknet_leaf_2_wb_clk_i _02760_ _00826_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14342_ _05123_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__nor2_1
X_11554_ _07377_ _07390_ _07458_ _07462_ _07464_ vssd1 vssd1 vccd1 vccd1 _07465_ sky130_fd_sc_hd__a2111o_4
XANTENNA__09290__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10505_ _06514_ _06517_ net382 vssd1 vssd1 vccd1 vccd1 _06518_ sky130_fd_sc_hd__o21a_2
X_17061_ clknet_leaf_175_wb_clk_i _02691_ _00757_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_14273_ _00034_ _00032_ _00031_ _04050_ vssd1 vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__nor4_1
X_11485_ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[16\] _07395_ net1003
+ vssd1 vssd1 vccd1 vccd1 _07396_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_150_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire587 _05756_ vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__clkbuf_1
X_16012_ net1114 vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__inv_2
X_13224_ net311 net2339 net350 vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10436_ net1019 _04922_ _04924_ net551 vssd1 vssd1 vccd1 vccd1 _06452_ sky130_fd_sc_hd__a211o_1
XFILLER_0_122_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08396__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13155_ net330 net2168 net445 vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12414__S net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10367_ _05841_ _05883_ _05881_ vssd1 vssd1 vccd1 vccd1 _06386_ sky130_fd_sc_hd__a21o_1
X_12106_ _07905_ _07906_ _07917_ _07910_ vssd1 vssd1 vccd1 vccd1 _07918_ sky130_fd_sc_hd__o31a_1
XANTENNA__11538__B _07447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10298_ _05899_ _06319_ vssd1 vssd1 vccd1 vccd1 _06320_ sky130_fd_sc_hd__nand2_4
X_13086_ _06655_ net2223 net454 vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__mux2_1
X_17963_ clknet_leaf_107_wb_clk_i net1961 _01659_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__dfrtp_1
X_12037_ _07842_ _07848_ _07450_ vssd1 vssd1 vccd1 vccd1 _07849_ sky130_fd_sc_hd__a21o_1
X_16914_ clknet_leaf_133_wb_clk_i _02544_ _00610_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_17894_ clknet_leaf_76_wb_clk_i _03237_ _01590_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13753__B _06387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16845_ clknet_leaf_159_wb_clk_i _02475_ _00541_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13245__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16776_ clknet_leaf_203_wb_clk_i _02406_ _00472_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13988_ net910 _03859_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[4\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15727_ net1292 vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12939_ net226 net2497 net469 vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_157_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08320__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15658_ net1245 vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_174_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14609_ net1216 vssd1 vssd1 vccd1 vccd1 _00239_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_174_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11207__A2 _07091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18377_ net1362 vssd1 vssd1 vccd1 vccd1 la_data_out[25] sky130_fd_sc_hd__buf_2
XANTENNA__08608__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09678__B net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15589_ net1249 vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__inv_2
XANTENNA__10415__A0 _06263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08130_ _04211_ _04216_ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17328_ clknet_leaf_137_wb_clk_i _02958_ _01024_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09820__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08061_ net1024 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__and2b_1
X_17259_ clknet_leaf_187_wb_clk_i _02889_ _00955_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09033__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10718__B2 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11729__A team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[10\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08963_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[15\]
+ net711 net695 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[15\]
+ _05025_ vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08894_ _04953_ _04955_ _04957_ _04959_ vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__or4_1
XFILLER_0_75_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10351__C1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout370_A net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13155__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout468_A net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09515_ net1017 net1014 net955 vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__o21a_1
X_18377__1362 vssd1 vssd1 vccd1 vccd1 _18377__1362/HI net1362 sky130_fd_sc_hd__conb_1
XFILLER_0_116_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12994__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout635_A _04313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09446_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[5\]
+ net817 net792 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10702__A2_N net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09377_ _05421_ vssd1 vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout802_A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout423_X net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08328_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[31\]
+ net772 _04409_ net855 vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09272__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10957__A1 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09811__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08259_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[31\]
+ net717 _04335_ _04341_ vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_62_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11270_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[98\] _07123_
+ _07130_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[98\] vssd1 vssd1
+ vccd1 vccd1 _07231_ sky130_fd_sc_hd__a22o_1
XANTENNA__09024__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout792_X net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08378__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10221_ net897 _06245_ _06246_ _06243_ vssd1 vssd1 vccd1 vccd1 _06247_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_37_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09754__D net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10152_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[29\] _06102_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[30\]
+ vssd1 vssd1 vccd1 vccd1 _06180_ sky130_fd_sc_hd__a21o_1
XANTENNA__09109__A _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10590__C1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09327__A1 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10083_ net891 _06108_ _06110_ net556 vssd1 vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__a211o_1
X_14960_ net1093 vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_54_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold9 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[8\]
+ vssd1 vssd1 vccd1 vccd1 net1423 sky130_fd_sc_hd__dlygate4sd3_1
X_13911_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[27\]
+ net559 net575 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[27\]
+ net986 vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__a221o_1
XANTENNA_input29_A DAT_I[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14891_ net1070 vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__inv_2
XANTENNA__13065__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16630_ clknet_leaf_150_wb_clk_i _02260_ _00326_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13842_ net1538 net579 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[20\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_69_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16561_ clknet_leaf_168_wb_clk_i _02191_ _00257_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13773_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[13\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[12\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[15\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__or4_1
XANTENNA__12634__A1 _07798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08838__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10985_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[15\] net564 _06964_
+ _06965_ vssd1 vssd1 vccd1 vccd1 _03421_ sky130_fd_sc_hd__a22o_1
X_15512_ net1161 vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__inv_2
X_18300_ net1392 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
XANTENNA__10645__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12724_ net306 net1971 net499 vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__mux2_1
X_16492_ clknet_leaf_1_wb_clk_i _02122_ _00188_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08683__A net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18231_ clknet_leaf_50_wb_clk_i net1489 _01926_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_15443_ net1258 vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__inv_2
X_12655_ net1921 _03691_ _03685_ vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__o21a_1
XANTENNA__12409__S net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18162_ clknet_leaf_152_wb_clk_i _03465_ _01858_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11606_ net1955 net1008 net344 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[19\]
+ vssd1 vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__a22o_1
X_15374_ net1190 vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__inv_2
X_12586_ net1834 _07793_ _03680_ vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09263__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10437__B _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17113_ clknet_leaf_9_wb_clk_i _02743_ _00809_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14325_ _05801_ _05768_ _05732_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__o2bb2a_1
X_18093_ clknet_leaf_66_wb_clk_i _03416_ _01789_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[10\]
+ sky130_fd_sc_hd__dfrtp_2
X_11537_ _07379_ _07447_ vssd1 vssd1 vccd1 vccd1 _07448_ sky130_fd_sc_hd__nor2_2
XFILLER_0_53_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire373 _05550_ vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__buf_4
Xhold409 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[61\] vssd1 vssd1
+ vccd1 vccd1 net1823 sky130_fd_sc_hd__dlygate4sd3_1
X_17044_ clknet_leaf_120_wb_clk_i _02674_ _00740_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_14256_ _00028_ _00039_ _04040_ vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09015__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13748__B _06481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11468_ _07369_ _07378_ vssd1 vssd1 vccd1 vccd1 _07379_ sky130_fd_sc_hd__nor2_4
XFILLER_0_111_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11549__A _07414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08369__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13207_ _06461_ net2538 net351 vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10419_ net337 _06253_ _06432_ net348 _06435_ vssd1 vssd1 vccd1 vccd1 _06436_ sky130_fd_sc_hd__o221a_1
X_14187_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[1\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[0\]
+ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[2\] vssd1 vssd1
+ vccd1 vccd1 _03996_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12570__A0 _03666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11399_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[15\] _07329_
+ vssd1 vssd1 vccd1 vccd1 _07330_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13138_ net247 net2198 net445 vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__mux2_1
XANTENNA__14311__A1 _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17946_ clknet_leaf_35_wb_clk_i _03285_ _01642_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13069_ net237 net2405 net454 vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__mux2_1
XANTENNA__14311__B2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[21\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1109 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2523 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10599__S net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09680__C net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08210__X _04293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17877_ clknet_leaf_91_wb_clk_i _03220_ _01573_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10333__C1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08541__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16828_ clknet_leaf_154_wb_clk_i _02458_ _00524_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_16759_ clknet_leaf_144_wb_clk_i _02389_ _00455_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09300_ _05334_ _05337_ _05338_ _05348_ vssd1 vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__or4_1
XFILLER_0_158_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09231_ _05281_ vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09162_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[11\]
+ net818 net774 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08113_ net1032 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__and2b_1
XFILLER_0_16_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09093_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[12\]
+ net682 net629 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[12\]
+ _05149_ vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout216_A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08044_ team_05_WB.instance_to_wrap.BUSY_O vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__inv_2
XANTENNA__09006__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold910 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2324 sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 net2335 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold932 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2346 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12010__C1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold943 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2357 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold954 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2368 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12561__A0 _03645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold965 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2379 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09574__D net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold976 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net2390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 net2401 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold998 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net2412 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12989__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09995_ _06020_ _06023_ net513 vssd1 vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_134_Left_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08780__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08946_ _04996_ _04997_ _05008_ _05009_ vssd1 vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__or4_1
XANTENNA__08768__A _04818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08877_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[17\]
+ net716 _04939_ _04943_ vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__o22a_2
XTAP_TAPCELL_ROW_4_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout752_A net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12577__X _03680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout540_X net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout638_X net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13613__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10770_ net2100 net305 net542 vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__mux2_1
XANTENNA__09493__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_143_Left_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14369__A1 _04128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09429_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[5\]
+ net670 net646 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[5\]
+ _05471_ vssd1 vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__a221o_1
XANTENNA__10097__X _06125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout805_X net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09749__D net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12440_ net919 _07860_ _07863_ _03659_ vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__and4_4
XANTENNA__09245__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08599__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12371_ net1737 _03651_ net216 vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14110_ _03971_ _03974_ vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__xor2_1
XFILLER_0_22_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11322_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[8\] _07101_ _07110_
+ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[48\] _07280_ vssd1 vssd1
+ vccd1 vccd1 _07281_ sky130_fd_sc_hd__a221o_1
XFILLER_0_22_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15090_ net1232 vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14041_ net910 _03910_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[6\]
+ sky130_fd_sc_hd__nor2_1
X_11253_ _07058_ _07085_ _07118_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[67\]
+ _07031_ vssd1 vssd1 vccd1 vccd1 _07215_ sky130_fd_sc_hd__a221o_1
XFILLER_0_127_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_152_Left_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10204_ _06151_ _06169_ net520 vssd1 vssd1 vccd1 vccd1 _06230_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11184_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[38\] _07097_
+ _07108_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[94\] vssd1 vssd1
+ vccd1 vccd1 _07149_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_128_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12899__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17800_ clknet_leaf_90_wb_clk_i _03143_ _01496_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[110\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_73_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10560__X _06570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10135_ _04470_ net510 net336 _06161_ _06162_ vssd1 vssd1 vccd1 vccd1 _06163_ sky130_fd_sc_hd__o221a_1
XANTENNA__08771__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15992_ net1128 vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_145_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17731_ clknet_leaf_86_wb_clk_i _03074_ _01427_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[41\]
+ sky130_fd_sc_hd__dfrtp_1
X_10066_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[17\] _06094_ vssd1
+ vssd1 vccd1 vccd1 _06095_ sky130_fd_sc_hd__and2_1
X_14943_ net1181 vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08523__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17662_ clknet_leaf_84_wb_clk_i _03005_ _01358_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[100\]
+ sky130_fd_sc_hd__dfrtp_1
X_14874_ net1062 vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_141_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16613_ clknet_leaf_19_wb_clk_i _02243_ _00309_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13825_ net1493 net578 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[3\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_173_1082 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17593_ clknet_leaf_73_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[30\]
+ _01289_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12928__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_161_Left_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13523__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10618__B1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16544_ clknet_leaf_126_wb_clk_i _02174_ _00240_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13756_ net922 _06320_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[24\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10968_ _06445_ _06951_ net956 vssd1 vssd1 vccd1 vccd1 _06952_ sky130_fd_sc_hd__mux2_1
XANTENNA__09484__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17499__Q team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12707_ net260 net2823 net496 vssd1 vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__mux2_1
XANTENNA__09302__A _05350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11291__B1 _07127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16475_ clknet_leaf_193_wb_clk_i _02105_ _00171_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13687_ net2238 net310 net384 vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10899_ net1044 _06181_ _06894_ net957 vssd1 vssd1 vccd1 vccd1 _06895_ sky130_fd_sc_hd__o211a_1
X_18214_ clknet_leaf_57_wb_clk_i net1461 _01909_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_15426_ net1128 vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__inv_2
X_12638_ _03666_ net1867 net201 vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09236__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15357_ net1087 vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__inv_2
X_18145_ clknet_leaf_17_wb_clk_i _03448_ _01841_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12569_ _03665_ net1871 net207 vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11594__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12791__A0 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11594__B2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[30\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14308_ _04071_ _04075_ _04076_ _04080_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__or4_1
X_18076_ clknet_leaf_84_wb_clk_i _00017_ _01772_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold206 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[123\] vssd1 vssd1
+ vccd1 vccd1 net1620 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_117_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08205__X _04288_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15288_ net1210 vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold217 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[13\] vssd1 vssd1
+ vccd1 vccd1 net1631 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09675__C net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold228 team_05_WB.instance_to_wrap.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 net1642
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_170_Left_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09539__A1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17027_ clknet_leaf_199_wb_clk_i _02657_ _00723_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_169_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14239_ net2665 _04021_ vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__nor2_1
Xhold239 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[21\] vssd1 vssd1
+ vccd1 vccd1 net1653 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_169_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18376__1361 vssd1 vssd1 vccd1 vccd1 _18376__1361/HI net1361 sky130_fd_sc_hd__conb_1
XFILLER_0_111_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout708 net710 vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout719 _04285_ vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_165_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[19\]
+ net837 net752 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08762__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12602__S net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09780_ _05442_ _05463_ vssd1 vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08731_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[21\]
+ net708 net630 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__a22o_1
X_17929_ clknet_leaf_43_wb_clk_i _03268_ _01625_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11726__B _07447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1290 net1291 vssd1 vssd1 vccd1 vccd1 net1290 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_89_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08662_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[23\]
+ net717 _04729_ _04735_ vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_89_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08593_ _04663_ _04665_ _04667_ _04668_ vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__or4_1
XANTENNA__13433__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15214__A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09475__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11282__B1 _07127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09569__D net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1083 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09214_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[10\]
+ net845 net809 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[10\]
+ _05265_ vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__a221o_1
XFILLER_0_134_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09145_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[11\]
+ net672 net617 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout500_A _07857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16045__A net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1242_A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09076_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[13\]
+ net821 net809 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[13\]
+ _05133_ vssd1 vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__a221o_1
XANTENNA__10364__Y _06384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09585__C net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08027_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[22\] vssd1
+ vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10093__A _05596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold740 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[15\] vssd1
+ vssd1 vccd1 vccd1 net2154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2165 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold762 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 net2176 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold773 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold784 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2198 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout490_X net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold795 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 net2209 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout967_A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_89_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13608__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08753__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12512__S net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09978_ net523 net362 vssd1 vssd1 vccd1 vccd1 _06007_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_51_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10560__A2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_18_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08929_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[16\]
+ net810 net771 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout755_X net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1440 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 net2854 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08505__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1451 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2865 sky130_fd_sc_hd__dlygate4sd3_1
X_11940_ net549 _07751_ vssd1 vssd1 vccd1 vccd1 _07752_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1462 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net2876 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1473 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2887 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1484 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2898 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1495 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2909 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout922_X net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11871_ _07648_ _07682_ vssd1 vssd1 vccd1 vccd1 _07683_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13343__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13610_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[14\]
+ net276 net395 vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__mux2_1
X_10822_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[11\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06819_ sky130_fd_sc_hd__nor2_1
X_14590_ net1054 vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11273__B1 _07129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13541_ net2751 net262 net401 vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__mux2_1
X_10753_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[1\] net904 _04247_
+ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[1\] vssd1 vssd1 vccd1
+ vccd1 _06752_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10268__A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16260_ net1116 vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13472_ net253 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[20\]
+ net408 vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__mux2_1
XANTENNA__09218__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10684_ _04173_ net902 net897 _06686_ _06684_ vssd1 vssd1 vccd1 vccd1 _06687_ sky130_fd_sc_hd__o221a_2
XFILLER_0_35_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15211_ net1070 vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__inv_2
X_12423_ net1688 _07812_ _03667_ vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__mux2_1
X_16191_ net1145 vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__inv_2
XFILLER_0_164_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15142_ net1231 vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__inv_2
X_12354_ _07993_ _03511_ vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11305_ _07254_ _07259_ _07260_ _07264_ vssd1 vssd1 vccd1 vccd1 _07265_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_75_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15073_ net1225 vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12285_ _03579_ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14024_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[15\] _04159_ vssd1
+ vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_147_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09792__A _05208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11236_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[36\] _07120_
+ _07197_ _07198_ vssd1 vssd1 vccd1 vccd1 _07199_ sky130_fd_sc_hd__a211o_1
XFILLER_0_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_123_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13518__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08744__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12422__S net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11167_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[15\] _07105_
+ _07110_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[55\] _07132_
+ vssd1 vssd1 vccd1 vccd1 _07133_ sky130_fd_sc_hd__a221o_1
XANTENNA__14278__B1 _06907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10118_ _05034_ net365 vssd1 vssd1 vccd1 vccd1 _06146_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11098_ _07046_ _07064_ vssd1 vssd1 vccd1 vccd1 _07065_ sky130_fd_sc_hd__and2_1
X_15975_ net1292 vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__inv_2
XANTENNA__10450__B _06464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17714_ clknet_leaf_92_wb_clk_i _03057_ _01410_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[88\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14926_ net1190 vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__inv_2
X_10049_ net379 net367 vssd1 vssd1 vccd1 vccd1 _06078_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_160_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11674__D_N net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13761__B _06185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17645_ clknet_leaf_69_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[12\]
+ _01341_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_14857_ net1222 vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_58_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13253__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13808_ net1611 net969 net724 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[19\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17576_ clknet_leaf_72_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[13\]
+ _01272_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_14788_ net1227 vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__inv_2
XANTENNA__09457__B1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13739_ net922 _06641_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[7\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16527_ clknet_leaf_138_wb_clk_i _02157_ _00223_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09209__B1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16458_ clknet_leaf_2_wb_clk_i _02088_ _00154_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15409_ net1132 vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__inv_2
X_16389_ clknet_leaf_180_wb_clk_i _02019_ _00085_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11567__A1 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11501__S net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12764__A0 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_162_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_84_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18128_ clknet_leaf_48_wb_clk_i _00024_ _01824_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08432__A1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10625__B _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18059_ net1037 _03397_ _01755_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_09901_ net377 _04878_ vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout505 net507 vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13428__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout516 net517 vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08735__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09393__C1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09832_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[20\]
+ net829 net748 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[20\]
+ _05861_ vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__a221o_1
Xfanout527 _05633_ vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_171_Right_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout538 _04276_ vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__buf_2
XANTENNA__10542__A2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout549 _07448_ vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__clkbuf_4
X_09763_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[0\]
+ net686 _05781_ _05783_ _05786_ vssd1 vssd1 vccd1 vccd1 _05794_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_77_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08714_ _04780_ _04782_ _04784_ _04786_ vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__or4_1
X_09694_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[1\]
+ net648 _05726_ net720 vssd1 vssd1 vccd1 vccd1 _05727_ sky130_fd_sc_hd__a211o_1
X_08645_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[23\]
+ net680 net630 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout450_A _03714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13163__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08576_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[25\]
+ net622 net604 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[25\]
+ _04651_ vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__a221o_1
XANTENNA__09448__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11255__B1 _07115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_136_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_136_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout715_A _04286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1078_X net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12507__S net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09128_ _05169_ _05171_ _05182_ _05183_ vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__or4_1
XFILLER_0_60_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09620__B1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09059_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[13\]
+ net617 _05117_ net720 vssd1 vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__a211o_1
XFILLER_0_20_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_92_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12070_ _07866_ _07869_ _07874_ vssd1 vssd1 vccd1 vccd1 _07882_ sky130_fd_sc_hd__and3_1
Xhold570 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1984 sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net1995 sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net2006 sky130_fd_sc_hd__dlygate4sd3_1
X_11021_ _06994_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[8\] net568
+ vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__mux2_1
XANTENNA__13338__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15760_ net1275 vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__inv_2
X_12972_ net228 net2229 net467 vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__mux2_1
XANTENNA__09687__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1270 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net2684 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input11_A DAT_I[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09151__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14711_ net1101 vssd1 vssd1 vccd1 vccd1 _00341_ sky130_fd_sc_hd__inv_2
Xhold1281 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2695 sky130_fd_sc_hd__dlygate4sd3_1
X_11923_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[2\] net997 vssd1
+ vssd1 vccd1 vccd1 _07735_ sky130_fd_sc_hd__nand2_2
X_15691_ net1160 vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__inv_2
Xhold1292 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net2706 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13073__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17430_ clknet_leaf_59_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[30\]
+ _01126_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14642_ net1238 vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__inv_2
X_11854_ _07628_ _07636_ _07632_ vssd1 vssd1 vccd1 vccd1 _07666_ sky130_fd_sc_hd__a21o_1
X_18375__1360 vssd1 vssd1 vccd1 vccd1 _18375__1360/HI net1360 sky130_fd_sc_hd__conb_1
XANTENNA__11246__B1 _07105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10805_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[18\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06802_ sky130_fd_sc_hd__nand2_1
X_17361_ clknet_leaf_36_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[25\]
+ _01057_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_14573_ net1079 vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11785_ _07576_ _07596_ _07559_ vssd1 vssd1 vccd1 vccd1 _07597_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_99_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12994__A0 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09787__A net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16312_ net1125 vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__inv_2
X_13524_ net2829 net326 net404 vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10736_ _04172_ net899 net895 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[2\]
+ _06735_ vssd1 vssd1 vccd1 vccd1 _06736_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_24_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17292_ clknet_leaf_0_wb_clk_i _02922_ _00988_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16243_ net1146 vssd1 vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__inv_2
X_13455_ net2011 net328 net414 vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12417__S net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10667_ _06668_ _06670_ _04264_ vssd1 vssd1 vccd1 vccd1 _06671_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_24_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12746__A0 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12406_ net500 net1748 net215 vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__mux2_1
X_16174_ net1153 vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_114_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13386_ net2444 net302 net421 vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10598_ net382 _06605_ vssd1 vssd1 vccd1 vccd1 _06606_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10221__A1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15125_ net1059 vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__inv_2
X_12337_ _03608_ _03631_ vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__or2_2
XANTENNA__12363__D _03657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08965__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__buf_2
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__buf_2
XFILLER_0_50_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15056_ net1182 vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13756__B _06320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12268_ _03561_ _03562_ vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__nand2_1
XANTENNA__13171__A0 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12660__B net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14007_ _03876_ _03877_ vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__nand2_1
XANTENNA__13248__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08717__A2 _04366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11219_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[45\] _07113_
+ _07118_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[69\] vssd1 vssd1
+ vccd1 vccd1 _07183_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_162_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09259__A1_N team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[21\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12199_ _07994_ _07998_ vssd1 vssd1 vccd1 vccd1 _08011_ sky130_fd_sc_hd__nor2_1
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__clkbuf_4
XANTENNA__09672__D net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09390__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire349_A _05305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11707__D _07478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15958_ net1272 vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__inv_2
XANTENNA__09142__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14909_ net1088 vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__inv_2
X_15889_ net1275 vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__inv_2
XANTENNA__12388__A _07478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08350__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08430_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[29\]
+ net593 _04503_ _04509_ vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__o22ai_4
X_17628_ clknet_leaf_59_wb_clk_i _02999_ _01324_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13226__A1 _06736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11237__B1 _07117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08361_ _04436_ _04438_ _04440_ _04441_ vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__or4_1
X_17559_ clknet_leaf_59_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[30\]
+ _01255_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08292_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[23\] _04149_
+ vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11488__A_N _07396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08956__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout302 _06655_ vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13158__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout498_A net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08708__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout313 net314 vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__clkbuf_2
Xfanout324 net325 vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__clkbuf_2
Xfanout335 _06065_ vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09582__D net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout346 _07473_ vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__clkbuf_4
Xfanout357 net358 vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__buf_2
XANTENNA_input3_A DAT_I[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09815_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[20\]
+ net660 net610 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__a22o_1
XANTENNA__09381__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12997__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout368 _05769_ vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout665_A _04305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09746_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[0\]
+ net881 _04287_ net859 vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__and4_1
XANTENNA__09669__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18340__1329 vssd1 vssd1 vccd1 vccd1 _18340__1329/HI net1329 sky130_fd_sc_hd__conb_1
XFILLER_0_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09677_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[1\]
+ net876 net869 net867 vssd1 vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__and4_1
XFILLER_0_55_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout453_X net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08341__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08628_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[24\]
+ net816 net792 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11228__B1 _07130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08559_ _04613_ _04632_ vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout620_X net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout718_X net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13621__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11570_ net1908 net1004 net727 _07438_ vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09841__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10521_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[14\] _06092_ vssd1
+ vssd1 vccd1 vccd1 _06533_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10451__A1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09757__D net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13240_ net247 net2645 net438 vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10452_ _06035_ _06037_ vssd1 vssd1 vccd1 vccd1 _06467_ sky130_fd_sc_hd__nand2_1
XFILLER_0_161_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08947__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13171_ net249 net2416 net442 vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__mux2_1
X_10383_ net896 _06401_ vssd1 vssd1 vccd1 vccd1 _06402_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12122_ _07927_ _07929_ _07923_ vssd1 vssd1 vccd1 vccd1 _07934_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_33_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_input59_A wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13068__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12053_ net547 _07541_ vssd1 vssd1 vccd1 vccd1 _07865_ sky130_fd_sc_hd__and2_1
X_16930_ clknet_leaf_5_wb_clk_i _02560_ _00626_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12900__A0 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11004_ net1045 _06979_ _06980_ vssd1 vssd1 vccd1 vccd1 _06981_ sky130_fd_sc_hd__a21bo_1
X_16861_ clknet_leaf_110_wb_clk_i _02491_ _00557_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_1071 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout880 net882 vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__clkbuf_2
X_15812_ net1300 vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__inv_2
Xfanout891 _04280_ vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12700__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16792_ clknet_leaf_28_wb_clk_i _02422_ _00488_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_15743_ net1292 vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__inv_2
X_12955_ net320 net2130 net469 vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11906_ net343 _07641_ _07679_ vssd1 vssd1 vccd1 vccd1 _07718_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_29_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15674_ net1261 vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__inv_2
X_12886_ net302 net2243 net477 vssd1 vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11219__B1 _07118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17413_ clknet_leaf_60_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[13\]
+ _01109_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_138_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10690__A1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14625_ net1236 vssd1 vssd1 vccd1 vccd1 _00255_ sky130_fd_sc_hd__inv_2
X_11837_ _07647_ _07644_ vssd1 vssd1 vccd1 vccd1 _07649_ sky130_fd_sc_hd__nand2b_1
X_18393_ net915 vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13531__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17344_ clknet_leaf_40_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[8\]
+ _01040_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14556_ net1083 vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_155_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ _07562_ _07579_ _07577_ vssd1 vssd1 vccd1 vccd1 _07580_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09832__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10719_ _06717_ _06719_ net382 vssd1 vssd1 vccd1 vccd1 _06720_ sky130_fd_sc_hd__o21a_2
X_13507_ net2062 net264 net404 vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17275_ clknet_leaf_190_wb_clk_i _02905_ _00971_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_14487_ net1101 vssd1 vssd1 vccd1 vccd1 _00117_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11699_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[20\] team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[24\]
+ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[27\] net993 vssd1 vssd1
+ vccd1 vccd1 _07511_ sky130_fd_sc_hd__o31a_1
XFILLER_0_141_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10993__A2 _06768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13438_ net2180 net246 net414 vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__mux2_1
X_16226_ net1205 vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08399__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16157_ net1166 vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08938__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13369_ net2047 net236 net421 vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15108_ net1230 vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__inv_2
X_16088_ net1308 vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__inv_2
XANTENNA__08213__X _04296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15039_ net1181 vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09363__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08299__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11170__A2 _07116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08571__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09600_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[2\]
+ net716 vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12610__S net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09531_ _05565_ _05566_ _05567_ _05568_ vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__or4_2
XANTENNA__09115__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08323__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09462_ _05489_ _05493_ _05501_ _05503_ vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__or4_1
XFILLER_0_149_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08413_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[29\]
+ _04417_ net744 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09393_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[6\]
+ net664 _05437_ net719 vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__a211o_1
XFILLER_0_19_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout246_A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13441__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08344_ net570 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__nor2_1
XANTENNA__09823__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08275_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[18\] _04357_
+ vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout413_A _03727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09577__D net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10984__A2 _06500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08929__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout201_X net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10736__A2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11468__Y _07379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout782_A net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1108 net1313 vssd1 vssd1 vccd1 vccd1 net1108 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1119 net1120 vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__buf_2
XFILLER_0_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout570_X net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08562__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout668_X net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13616__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11925__A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12520__S net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout198 net200 vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09106__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09729_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[0\]
+ net738 _05738_ _05743_ _05750_ vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__13989__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_151_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_151_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout835_X net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12740_ net258 net2359 net492 vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10672__A1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12671_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[18\]
+ net339 vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14410_ net953 _04360_ _04346_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[23\]
+ sky130_fd_sc_hd__a21o_1
XANTENNA__13351__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11622_ net138 net1008 net344 net2012 vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15390_ net1073 vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09814__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14341_ _05596_ net533 net373 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__o2bb2a_1
X_11553_ _07348_ _07353_ _07434_ _07463_ vssd1 vssd1 vccd1 vccd1 _07464_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_133_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10424__B2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[19\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire533 _05575_ vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__buf_4
XFILLER_0_107_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10504_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[15\] net903 net965
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[15\] _06516_ vssd1
+ vssd1 vccd1 vccd1 _06517_ sky130_fd_sc_hd__a221o_1
X_17060_ clknet_leaf_182_wb_clk_i _02690_ _00756_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_14272_ _04042_ _00037_ _00036_ _04049_ vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__or4_1
XFILLER_0_80_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11484_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[16\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[16\]
+ net1031 vssd1 vssd1 vccd1 vccd1 _07395_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_150_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16011_ net1114 vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_150_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13223_ net328 net2499 net352 vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire588 net589 vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13913__A2 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10435_ _06284_ _06450_ net370 vssd1 vssd1 vccd1 vccd1 _06451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09129__X team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[12\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09593__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13154_ net313 net2863 net446 vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10366_ net2003 net228 net541 vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_29_Left_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12105_ _07902_ _07908_ vssd1 vssd1 vccd1 vccd1 _07917_ sky130_fd_sc_hd__nor2_1
X_13085_ net295 net2632 net455 vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__mux2_1
X_17962_ clknet_leaf_108_wb_clk_i net2013 _01658_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__dfrtp_1
X_10297_ _05894_ _05898_ vssd1 vssd1 vccd1 vccd1 _06319_ sky130_fd_sc_hd__nand2_1
X_12036_ _07377_ _07846_ vssd1 vssd1 vccd1 vccd1 _07848_ sky130_fd_sc_hd__or2_1
X_16913_ clknet_leaf_168_wb_clk_i _02543_ _00609_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17893_ clknet_leaf_101_wb_clk_i _03236_ _01589_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_109_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08553__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12430__S _03668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16844_ clknet_leaf_0_wb_clk_i _02474_ _00540_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_16775_ clknet_leaf_203_wb_clk_i _02405_ _00471_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13987_ _03857_ _03858_ _03839_ vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_105_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15726_ net1256 vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__inv_2
X_12938_ net230 net2401 net470 vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_157_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_38_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10663__A1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_122_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15657_ net1249 vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12869_ net236 net2625 net477 vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13261__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14608_ net1092 vssd1 vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_174_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18376_ net1361 vssd1 vssd1 vccd1 vccd1 la_data_out[24] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_174_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15588_ net1249 vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__inv_2
XANTENNA__09678__C net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09040__A team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[14\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17327_ clknet_leaf_135_wb_clk_i _02957_ _01023_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11612__B1 _07472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08084__A2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[19\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14539_ net1077 vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08060_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[31\] net1027
+ net974 _04179_ vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__a22o_1
XANTENNA__09975__A _05731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17258_ clknet_leaf_195_wb_clk_i _02888_ _00954_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16209_ net1232 vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__inv_2
XANTENNA__13904__A2 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12605__S _03680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17189_ clknet_leaf_18_wb_clk_i _02819_ _00885_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_47_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09039__X team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[14\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08792__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08962_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[15\]
+ net682 net610 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__a22o_1
X_18354__1339 vssd1 vssd1 vccd1 vccd1 _18354__1339/HI net1339 sky130_fd_sc_hd__conb_1
XANTENNA__09336__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08893_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[17\]
+ net849 net752 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[17\]
+ _04958_ vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout196_A _06184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08544__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13436__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09514_ _05551_ _05552_ vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_56_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_918 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09445_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[5\]
+ net804 net743 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1272_A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13171__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout249_X net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09376_ net375 _05419_ vssd1 vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__and2_1
XFILLER_0_163_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08327_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[31\]
+ net769 net765 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11603__B1 _07472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout416_X net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10957__A2 _06408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08258_ _04337_ _04338_ _04339_ _04340_ vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__or4_1
XFILLER_0_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_65_Left_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12515__S _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08189_ _04267_ _04271_ vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__or2_2
XFILLER_0_43_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10220_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[28\] net903 net965
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[28\] vssd1 vssd1
+ vccd1 vccd1 _06246_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_123_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout785_X net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10151_ _06003_ _06141_ _06178_ _06111_ vssd1 vssd1 vccd1 vccd1 _06179_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_37_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09327__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13854__B net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10082_ net891 _06109_ vssd1 vssd1 vccd1 vccd1 _06110_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_54_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13346__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13910_ net1812 net982 _03791_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[26\]
+ sky130_fd_sc_hd__o21a_1
X_14890_ net1121 vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11374__B net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13841_ net1502 net579 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[19\]
+ sky130_fd_sc_hd__and2_1
X_13772_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[9\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[8\] team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[11\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__or4_1
X_16560_ clknet_leaf_123_wb_clk_i _02190_ _00256_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10984_ net960 _06500_ net565 vssd1 vssd1 vccd1 vccd1 _06965_ sky130_fd_sc_hd__a21oi_1
X_15511_ net1167 vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__inv_2
XANTENNA__10645__A1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12723_ net326 net1915 net499 vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16491_ clknet_leaf_187_wb_clk_i _02121_ _00187_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13081__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18230_ clknet_leaf_52_wb_clk_i net1494 _01925_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_15442_ net1259 vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__inv_2
X_12654_ _07346_ _03686_ vssd1 vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12398__A1 _07821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_152_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11605_ net1840 net1009 net344 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18161_ clknet_leaf_124_wb_clk_i _03464_ _01857_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_12585_ _03657_ net1894 net204 vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15373_ net1088 vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17112_ clknet_leaf_28_wb_clk_i _02742_ _00808_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11536_ _07377_ _07390_ _07420_ _07446_ vssd1 vssd1 vccd1 vccd1 _07447_ sky130_fd_sc_hd__a211o_4
XFILLER_0_81_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14324_ _05442_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[6\]
+ net374 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[5\] vssd1
+ vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__o22a_1
X_18092_ clknet_leaf_66_wb_clk_i _03415_ _01788_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_29_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13347__A0 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwire374 _05483_ vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__clkbuf_4
X_14255_ _00027_ _00026_ _00025_ _04039_ vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__or4_1
X_17043_ clknet_leaf_166_wb_clk_i _02673_ _00739_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11467_ _07377_ _07363_ vssd1 vssd1 vccd1 vccd1 _07378_ sky130_fd_sc_hd__nand2b_2
XANTENNA__12425__S net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10293__X _06316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13206_ net255 net2338 net350 vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10418_ net334 _06255_ _06355_ _06252_ _06434_ vssd1 vssd1 vccd1 vccd1 _06435_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_78_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14186_ _07026_ net728 _03995_ vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__and3_1
XANTENNA__11549__B _07438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11398_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[14\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[13\]
+ _07328_ vssd1 vssd1 vccd1 vccd1 _07329_ sky130_fd_sc_hd__and3_1
XANTENNA__11373__A2 _06769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08774__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13137_ net228 net2481 net446 vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__mux2_1
X_10349_ _05890_ _05982_ vssd1 vssd1 vccd1 vccd1 _06369_ sky130_fd_sc_hd__xnor2_4
XANTENNA__09318__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17945_ clknet_leaf_35_wb_clk_i _03284_ _01641_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13068_ net240 net2318 net454 vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__mux2_1
XANTENNA__14311__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[22\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08526__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13256__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12019_ _07822_ _07824_ _07829_ _07830_ vssd1 vssd1 vccd1 vccd1 _07831_ sky130_fd_sc_hd__and4b_1
XFILLER_0_174_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17876_ clknet_leaf_88_wb_clk_i _03219_ _01572_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_79_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_136_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09680__D net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16827_ clknet_leaf_192_wb_clk_i _02457_ _00523_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10396__A1_N _05881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16758_ clknet_leaf_138_wb_clk_i _02388_ _00454_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15709_ net1165 vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__inv_2
X_16689_ clknet_leaf_122_wb_clk_i _02319_ _00385_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11504__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09230_ _05280_ _05256_ vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_61_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10187__Y _06214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12389__A1 _03664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09161_ _05215_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[11\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_56_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18359_ net1344 vssd1 vssd1 vccd1 vccd1 la_data_out[7] sky130_fd_sc_hd__buf_2
XFILLER_0_43_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08112_ net1028 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[5\]
+ net975 _04205_ vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09092_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[12\]
+ net704 net652 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_831 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08043_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[4\] vssd1
+ vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold900 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 net2314 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold911 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2325 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout209_A _03676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold922 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net2336 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12010__B1 _07774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09557__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold933 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net2347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold944 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold955 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 net2369 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10167__A3 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold966 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net2391 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1020_A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold988 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net2402 sky130_fd_sc_hd__dlygate4sd3_1
X_09994_ _06021_ _06022_ vssd1 vssd1 vccd1 vccd1 _06023_ sky130_fd_sc_hd__nand2_1
Xhold999 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net2413 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09309__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08945_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[16\]
+ net774 net768 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[16\]
+ _04993_ vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__a221o_1
XANTENNA__10650__Y _06655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout480_A net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout578_A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13166__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08876_ _04930_ _04931_ _04941_ _04942_ vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__or4_1
XANTENNA__10324__B1 _04265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09190__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout745_A _04417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10627__A1 _06338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08296__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09428_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[5\]
+ net654 net604 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09359_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[7\]
+ net757 net742 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[7\]
+ _05404_ vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout700_X net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12370_ net1678 _03662_ net216 vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11321_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[32\] _07097_
+ _07102_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[104\] vssd1
+ vssd1 vccd1 vccd1 _07280_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14040_ _03883_ _03909_ vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__nand2_1
X_11252_ _07031_ _07085_ vssd1 vssd1 vccd1 vccd1 _07214_ sky130_fd_sc_hd__or2_1
XANTENNA__09548__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12552__A1 _07793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10203_ _06225_ _06228_ net370 vssd1 vssd1 vccd1 vccd1 _06229_ sky130_fd_sc_hd__mux2_1
XANTENNA__08756__B1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_113_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11183_ _07133_ _07134_ _07148_ _07090_ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_128_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input41_A wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10134_ net1020 _04468_ _04469_ net552 vssd1 vssd1 vccd1 vccd1 _06162_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_73_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15991_ net1128 vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__inv_2
XANTENNA__08508__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13076__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17730_ clknet_leaf_94_wb_clk_i _03073_ _01426_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_145_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10065_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[16\] team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[15\]
+ _06093_ vssd1 vssd1 vccd1 vccd1 _06094_ sky130_fd_sc_hd__and3_1
X_14942_ net1054 vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__inv_2
X_17661_ clknet_leaf_102_wb_clk_i _03004_ _01357_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[99\]
+ sky130_fd_sc_hd__dfrtp_1
X_14873_ net1057 vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__inv_2
XANTENNA_output128_A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16612_ clknet_leaf_182_wb_clk_i _02242_ _00308_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13824_ net1473 net581 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[2\]
+ sky130_fd_sc_hd__and2_1
X_17592_ clknet_leaf_113_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[29\]
+ _01288_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_173_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10618__A1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16543_ clknet_leaf_152_wb_clk_i _02173_ _00239_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13755_ _05212_ _06350_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[23\]
+ sky130_fd_sc_hd__and2_1
X_10967_ net1042 _06869_ _06949_ _06950_ vssd1 vssd1 vccd1 vccd1 _06951_ sky130_fd_sc_hd__a31o_1
XFILLER_0_85_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12706_ net265 net2260 net496 vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16474_ clknet_leaf_12_wb_clk_i _02104_ _00170_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10898_ net1044 _06886_ _06893_ vssd1 vssd1 vccd1 vccd1 _06894_ sky130_fd_sc_hd__nand3_1
XFILLER_0_127_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13686_ net2039 net331 net385 vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__mux2_1
X_18213_ clknet_leaf_56_wb_clk_i net1821 _01908_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18353__1338 vssd1 vssd1 vccd1 vccd1 _18353__1338/HI net1338 sky130_fd_sc_hd__conb_1
X_15425_ net1123 vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12637_ _03665_ net1846 _03683_ vssd1 vssd1 vccd1 vccd1 _03008_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15320__A net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18144_ clknet_leaf_148_wb_clk_i _03447_ _01840_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12568_ _03605_ net1740 net206 vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__mux2_1
XANTENNA__13759__B _06907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_152_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15356_ net1064 vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12663__B net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11594__A2 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11519_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[24\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[24\]
+ net1033 vssd1 vssd1 vccd1 vccd1 _07430_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_152_Right_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14307_ _04072_ _04073_ _04074_ _04079_ vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__or4_1
X_18075_ clknet_leaf_85_wb_clk_i _00016_ _01771_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_145_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12499_ net1721 _03605_ net210 vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_117_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15287_ net1097 vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__inv_2
Xhold207 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[19\] vssd1 vssd1
+ vccd1 vccd1 net1621 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09675__D net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold218 net98 vssd1 vssd1 vccd1 vccd1 net1632 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold229 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[101\] vssd1 vssd1
+ vccd1 vccd1 net1643 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09539__A2 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17026_ clknet_leaf_4_wb_clk_i _02656_ _00722_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_14238_ net2000 _04022_ vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_169_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08747__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14169_ team_05_WB.instance_to_wrap.CPU_DAT_O\[18\] net504 net908 vssd1 vssd1 vccd1
+ vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[18\] sky130_fd_sc_hd__and3_1
XANTENNA__16151__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08211__A2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout709 net710 vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__buf_4
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08730_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[21\]
+ net661 net638 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[21\]
+ _04801_ vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__a221o_1
X_17928_ clknet_leaf_43_wb_clk_i _03267_ _01624_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09172__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1280 net1312 vssd1 vssd1 vccd1 vccd1 net1280 sky130_fd_sc_hd__buf_4
Xfanout1291 net1311 vssd1 vssd1 vccd1 vccd1 net1291 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_1_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08661_ _04731_ _04732_ _04733_ _04734_ vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__or4_1
X_17859_ clknet_leaf_77_wb_clk_i _03202_ _01555_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[41\]
+ sky130_fd_sc_hd__dfrtp_1
X_08592_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[25\]
+ net789 net765 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[25\]
+ _04657_ vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__a221o_1
XANTENNA__10609__B2 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_191_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09213_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[10\]
+ net801 net745 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout326_A net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09144_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[11\]
+ net668 net660 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[11\]
+ _05198_ vssd1 vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__a221o_1
XANTENNA__15230__A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08986__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09075_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[13\]
+ net815 net787 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__a22o_1
XFILLER_0_170_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09585__D net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08026_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[24\] vssd1
+ vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__inv_2
Xhold730 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold741 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2155 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08738__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout695_A net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold752 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 net2166 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold763 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2177 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold774 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 net2188 sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2199 sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net2210 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout483_X net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout862_A net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09977_ _05596_ net362 vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_51_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08928_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[28\] net966
+ net955 _04992_ _04345_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[16\]
+ sky130_fd_sc_hd__a221o_1
Xhold1430 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2844 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09163__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1441 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 net2855 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1452 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 net2866 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout650_X net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1463 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2877 sky130_fd_sc_hd__dlygate4sd3_1
X_08859_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[17\]
+ net671 net655 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__a22o_1
Xhold1474 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2888 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout748_X net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08910__B1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13624__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1485 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net2899 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_58_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11870_ _07681_ vssd1 vssd1 vccd1 vccd1 _07682_ sky130_fd_sc_hd__inv_2
Xhold1496 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net2910 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10821_ _06816_ _06817_ vssd1 vssd1 vccd1 vccd1 _06818_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout915_X net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13540_ net1954 net264 net400 vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__mux2_1
X_10752_ _06738_ _06750_ net536 vssd1 vssd1 vccd1 vccd1 _06751_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13471_ net247 net2767 net410 vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__mux2_1
X_10683_ _06087_ _06685_ vssd1 vssd1 vccd1 vccd1 _06686_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11025__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12422_ _03645_ net1889 net215 vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15210_ net1110 vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__inv_2
X_16190_ net1145 vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__inv_2
XANTENNA__08306__X _04388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08977__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12353_ _03643_ _03644_ _03645_ _03647_ vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__and4_1
X_15141_ net1193 vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08441__A2 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11304_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[49\] _07110_
+ _07250_ _07263_ vssd1 vssd1 vccd1 vccd1 _07264_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_75_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15072_ net1195 vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12284_ _08004_ _08006_ _03577_ vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_75_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12525__A1 _03632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14023_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[15\] _04159_ vssd1
+ vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08729__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11235_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[44\] _07113_
+ _07125_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[20\] _07031_
+ vssd1 vssd1 vccd1 vccd1 _07198_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_147_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12703__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11166_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[7\] _07100_ _07128_
+ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[71\] vssd1 vssd1 vccd1
+ vccd1 _07132_ sky130_fd_sc_hd__a22o_1
XANTENNA__14278__A1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10731__B net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10117_ _04989_ net364 vssd1 vssd1 vccd1 vccd1 _06145_ sky130_fd_sc_hd__or2_1
XANTENNA__10223__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11097_ _04161_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[1\]
+ _04164_ _07048_ _07054_ vssd1 vssd1 vccd1 vccd1 _07064_ sky130_fd_sc_hd__a41o_1
X_15974_ net1267 vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__inv_2
XANTENNA__09154__B1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[20\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17713_ clknet_leaf_98_wb_clk_i _03056_ _01409_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[87\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14925_ net1081 vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__inv_2
X_10048_ _04656_ net363 vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_160_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_4_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_160_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold90 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[24\]
+ vssd1 vssd1 vccd1 vccd1 net1504 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13534__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17644_ clknet_leaf_68_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[11\]
+ _01340_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_14856_ net1219 vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__inv_2
XANTENNA__12658__B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13807_ net1590 net972 net724 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[18\]
+ sky130_fd_sc_hd__and3_1
X_17575_ clknet_leaf_73_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[12\]
+ _01271_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14787_ net1207 vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__inv_2
X_11999_ _07809_ _07810_ _07799_ vssd1 vssd1 vccd1 vccd1 _07811_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_11_Left_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16526_ clknet_leaf_171_wb_clk_i _02156_ _00222_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13738_ net922 _06658_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[6\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_133_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_978 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16457_ clknet_leaf_20_wb_clk_i _02087_ _00153_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_119_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13669_ net2376 net246 net385 vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15408_ net1138 vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16388_ clknet_leaf_182_wb_clk_i _02018_ _00084_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09686__C net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08968__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18127_ clknet_leaf_48_wb_clk_i _00023_ _01823_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15339_ net1077 vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08432__A2 _04510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18058_ net1037 _03396_ _01754_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12516__A1 _03657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09900_ _04756_ _04758_ vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__nand2_4
XPHY_EDGE_ROW_20_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17009_ clknet_leaf_118_wb_clk_i _02639_ _00705_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12613__S net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10527__B1 _04279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout506 net507 vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09831_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[20\]
+ net849 net782 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__a22o_1
Xfanout517 net522 vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__buf_2
Xfanout528 net532 vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__clkbuf_4
Xfanout539 net542 vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__buf_6
XFILLER_0_158_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09762_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[0\]
+ net633 _05772_ _05776_ _05789_ vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09145__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08713_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[22\]
+ net780 net765 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[22\]
+ _04785_ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__a221o_1
X_09693_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[1\]
+ net703 net652 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__a22o_1
XANTENNA__14326__A2_N _05208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08499__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13444__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11753__A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08644_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[23\]
+ net684 net623 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08575_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[25\]
+ net685 net612 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout443_A _03716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1185_A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout610_A _04319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08671__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout708_A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_176_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_176_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08959__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09127_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[12\]
+ net798 net794 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[12\]
+ _05170_ vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_105_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_105_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09081__C1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09893__A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09058_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[13\]
+ net691 net637 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12507__A1 _03623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout698_X net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13619__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12523__S net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold560 team_05_WB.instance_to_wrap.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 net1974
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold571 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net1985 sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ net963 _06623_ _06993_ vssd1 vssd1 vccd1 vccd1 _06994_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09384__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold582 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net1996 sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2007 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_10__f_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18352__1337 vssd1 vssd1 vccd1 vccd1 _18352__1337/HI net1337 sky130_fd_sc_hd__conb_1
XANTENNA__09136__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12971_ net231 net2735 net467 vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__mux2_1
Xhold1260 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2674 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13354__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14710_ net1091 vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__inv_2
Xhold1271 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2685 sky130_fd_sc_hd__dlygate4sd3_1
X_11922_ _07691_ _07698_ vssd1 vssd1 vccd1 vccd1 _07734_ sky130_fd_sc_hd__xnor2_2
Xhold1282 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2696 sky130_fd_sc_hd__dlygate4sd3_1
X_15690_ net1166 vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__inv_2
Xhold1293 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2707 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14641_ net1192 vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11853_ _07628_ _07635_ vssd1 vssd1 vccd1 vccd1 _07665_ sky130_fd_sc_hd__xnor2_2
XANTENNA__10279__A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10804_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[19\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[19\]
+ vssd1 vssd1 vccd1 vccd1 _06801_ sky130_fd_sc_hd__and2_1
X_17360_ clknet_leaf_42_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[24\]
+ _01056_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14572_ net1070 vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__inv_2
X_11784_ _07594_ _07595_ _07580_ vssd1 vssd1 vccd1 vccd1 _07596_ sky130_fd_sc_hd__a21o_1
XFILLER_0_67_364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08972__A _05034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16311_ net1118 vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13523_ net1841 net322 net404 vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17291_ clknet_leaf_188_wb_clk_i _02921_ _00987_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10735_ _06731_ _06732_ _06734_ net538 vssd1 vssd1 vccd1 vccd1 _06735_ sky130_fd_sc_hd__a31o_1
XFILLER_0_138_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08662__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16242_ net1144 vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_136_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10666_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[6\] net906 net897
+ _06669_ vssd1 vssd1 vccd1 vccd1 _06670_ sky130_fd_sc_hd__o2bb2a_1
X_13454_ net2711 net315 net415 vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12405_ _07858_ _07863_ _03659_ vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__nand3b_4
XFILLER_0_3_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16173_ net1152 vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13385_ net2138 net294 net422 vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__mux2_1
X_10597_ _06601_ _06604_ vssd1 vssd1 vccd1 vccd1 _06605_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_114_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08414__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10757__B1 _06051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15124_ net1066 vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__inv_2
X_12336_ net544 _07475_ _03552_ vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__or3_1
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__buf_2
XANTENNA__13529__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12433__S _03667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12267_ _07970_ _03557_ _03554_ vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__a21bo_1
X_15055_ net1286 vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__inv_2
X_11218_ _07171_ _07173_ _07181_ vssd1 vssd1 vccd1 vccd1 _07182_ sky130_fd_sc_hd__or3_1
X_14006_ _03848_ _03875_ _03849_ vssd1 vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__or3b_1
X_12198_ _07987_ _08009_ _08007_ _08000_ vssd1 vssd1 vccd1 vccd1 _08010_ sky130_fd_sc_hd__a2bb2o_1
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_162_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__clkbuf_4
X_11149_ _07060_ _07114_ vssd1 vssd1 vccd1 vccd1 _07115_ sky130_fd_sc_hd__nor2_4
XANTENNA__09127__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15957_ net1269 vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__inv_2
XANTENNA__13264__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14908_ net1083 vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__inv_2
X_15888_ net1264 vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09043__A _05078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17627_ clknet_leaf_59_wb_clk_i _02998_ _01323_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14839_ net1096 vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13226__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12434__A0 _03650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08360_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[30\]
+ net713 net680 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[30\]
+ _04429_ vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__a221o_1
XANTENNA__09978__A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17558_ clknet_leaf_59_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[29\]
+ _01254_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08638__C1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_3_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16509_ clknet_leaf_128_wb_clk_i _02139_ _00205_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_08291_ net948 net1014 net933 vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__and3_4
XANTENNA__12608__S _03680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17489_ clknet_leaf_42_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[24\]
+ _01185_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08653__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09850__A1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08405__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_6__f_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13439__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout303 net304 vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__clkbuf_2
Xfanout314 net316 vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11173__B1 _07129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout325 net327 vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout393_A _03732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout336 _06065_ vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__buf_2
Xfanout347 _06508_ vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__buf_2
X_09814_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[20\]
+ net699 net602 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[20\]
+ _05844_ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__a221o_1
Xfanout358 _07469_ vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout369 _05577_ vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1100_A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09118__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09745_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[0\]
+ net880 net863 net859 vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout560_A net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13174__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout658_A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09676_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[1\]
+ net883 net864 net862 vssd1 vssd1 vccd1 vccd1 _05709_ sky130_fd_sc_hd__and4_1
XFILLER_0_55_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08166__D_N net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08627_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[24\]
+ net819 net779 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10099__A net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08892__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout446_X net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12425__A0 _03664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08558_ _04633_ vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10436__C1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12518__S _03676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08489_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[27\]
+ net673 net626 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[27\]
+ _04566_ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout613_X net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08644__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10520_ _06522_ _06530_ _06531_ net536 vssd1 vssd1 vccd1 vccd1 _06532_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10451_ net892 _06463_ _06465_ net554 vssd1 vssd1 vccd1 vccd1 _06466_ sky130_fd_sc_hd__a211o_1
XFILLER_0_162_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13170_ net227 net2652 net442 vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__mux2_1
X_10382_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[21\] _06097_ vssd1
+ vssd1 vccd1 vccd1 _06401_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_131_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12121_ _07927_ _07929_ _07923_ vssd1 vssd1 vccd1 vccd1 _07933_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13349__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09357__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12052_ net543 _07523_ vssd1 vssd1 vccd1 vccd1 _07864_ sky130_fd_sc_hd__or2_4
Xhold390 net91 vssd1 vssd1 vccd1 vccd1 net1804 sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ net1045 _06091_ _06586_ net959 vssd1 vssd1 vccd1 vccd1 _06980_ sky130_fd_sc_hd__o31a_1
Xclkbuf_leaf_73_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16860_ clknet_leaf_158_wb_clk_i _02490_ _00556_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10911__A0 _06219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout870 _04287_ vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__buf_2
XFILLER_0_99_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15811_ net1305 vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__inv_2
Xfanout881 net882 vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__buf_1
Xfanout892 _04279_ vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__clkbuf_4
X_16791_ clknet_leaf_144_wb_clk_i _02421_ _00487_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13084__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15742_ net1267 vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__inv_2
X_12954_ net302 net2920 net469 vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__mux2_1
Xhold1090 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2504 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11905_ _07716_ vssd1 vssd1 vccd1 vccd1 _07717_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_29_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15673_ net1261 vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12001__B _07475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12885_ net297 net2883 net478 vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__mux2_1
XANTENNA__08883__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17412_ clknet_leaf_60_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[12\]
+ _01108_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12416__A0 _03610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ net1198 vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__inv_2
X_18392_ net915 vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__clkbuf_1
X_11836_ _07644_ _07645_ _07647_ vssd1 vssd1 vccd1 vccd1 _07648_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_103_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ clknet_leaf_41_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[7\]
+ _01039_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14555_ net1099 vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__inv_2
XANTENNA__12428__S _03667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08635__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10737__A _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11767_ _07572_ _07578_ vssd1 vssd1 vccd1 vccd1 _07579_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_155_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13506_ net1986 net256 net405 vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__mux2_1
X_10718_ _04247_ _06085_ _06718_ net905 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06719_ sky130_fd_sc_hd__a32o_1
X_17274_ clknet_leaf_12_wb_clk_i _02904_ _00970_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_14486_ net1084 vssd1 vssd1 vccd1 vccd1 _00116_ sky130_fd_sc_hd__inv_2
X_11698_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[24\] net1000 vssd1
+ vssd1 vccd1 vccd1 _07510_ sky130_fd_sc_hd__and2_1
XFILLER_0_114_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16225_ net1204 vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13437_ net2035 net228 net414 vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10649_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[7\] net906 net897
+ _06653_ vssd1 vssd1 vccd1 vccd1 _06654_ sky130_fd_sc_hd__o2bb2a_1
X_16156_ net1253 vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13368_ net1992 net238 net421 vssd1 vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__mux2_1
XANTENNA__12671__B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09060__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15107_ net1197 vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__inv_2
XANTENNA__13259__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12319_ _03608_ _03613_ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__or2_4
X_16087_ net1308 vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__inv_2
XANTENNA__09683__D net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13299_ net2207 net218 net430 vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__mux2_1
XANTENNA__09348__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15038_ net1054 vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__inv_2
XANTENNA__14341__B1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16989_ clknet_leaf_108_wb_clk_i _02619_ _00685_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09530_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[3\]
+ net845 net833 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[3\]
+ _05558_ vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__a221o_1
XANTENNA__09520__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09461_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[5\]
+ net820 net735 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[5\]
+ _05502_ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__a221o_1
XANTENNA__10130__A1 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08874__A2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12407__A0 _03661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08412_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[29\]
+ net773 net733 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09392_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[6\]
+ net643 net601 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08343_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[31\]
+ net592 _04399_ _04424_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[31\]
+ sky130_fd_sc_hd__o22a_4
XFILLER_0_4_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13080__A0 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08626__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08274_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[17\] _04356_
+ vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_15_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11630__A1 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11630__B2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18351__1336 vssd1 vssd1 vccd1 vccd1 _18351__1336/HI net1336 sky130_fd_sc_hd__conb_1
XFILLER_0_46_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_918 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1050_A team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout406_A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09051__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13169__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09339__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout396_X net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout775_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1109 net1111 vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11697__A1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[19\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12801__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout199 net200 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11449__A1 _07346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09728_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[0\]
+ net846 _05746_ _05749_ _05752_ vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_96_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout730_X net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09659_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[1\]
+ net798 net782 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[1\]
+ _05687_ vssd1 vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__a221o_1
XANTENNA__08865__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13632__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout828_X net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12670_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[19\]
+ net339 vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_191_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_191_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11621_ net1960 net1008 net345 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[9\]
+ vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_61_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_120_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_120_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_108_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08617__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10424__A2 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14340_ _05208_ net535 _05256_ net534 vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__o22a_1
X_11552_ _07357_ _07360_ _07431_ _07436_ vssd1 vssd1 vccd1 vccd1 _07463_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_133_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08027__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[22\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09290__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire523 _05666_ vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__buf_2
X_10503_ net896 _06515_ vssd1 vssd1 vccd1 vccd1 _06516_ sky130_fd_sc_hd__nor2_1
Xwire534 _05279_ vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__buf_4
X_14271_ team_05_WB.instance_to_wrap.total_design.key_confirm _00035_ _00033_ _04217_
+ vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__or4b_1
X_11483_ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[25\] _07393_ net1001
+ vssd1 vssd1 vccd1 vccd1 _07394_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_150_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16010_ net1114 vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__inv_2
XANTENNA_input71_A wbs_cyc_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13222_ _06687_ net353 _03719_ vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__o21ai_1
X_10434_ _06377_ _06448_ net530 vssd1 vssd1 vccd1 vccd1 _06450_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_150_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire589 _05694_ vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10563__Y _06572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13079__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13153_ net319 net2428 net445 vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__mux2_1
XANTENNA__08250__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10365_ net383 _06384_ vssd1 vssd1 vccd1 vccd1 _06385_ sky130_fd_sc_hd__and2_1
XANTENNA__10292__A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_5__f_wb_clk_i_X clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12104_ _07914_ _07913_ _07912_ vssd1 vssd1 vccd1 vccd1 _07916_ sky130_fd_sc_hd__nand3b_2
XANTENNA__14323__B1 _05442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13084_ net300 net2535 net454 vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__mux2_1
X_17961_ clknet_leaf_108_wb_clk_i net1931 _01657_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__dfrtp_1
X_10296_ net2320 net240 net541 vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12035_ _07377_ _07450_ _07845_ _07369_ vssd1 vssd1 vccd1 vccd1 _07847_ sky130_fd_sc_hd__or4b_2
X_16912_ clknet_leaf_167_wb_clk_i _02542_ _00608_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_17892_ clknet_leaf_88_wb_clk_i _03235_ _01588_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12711__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_69_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16843_ clknet_leaf_186_wb_clk_i _02473_ _00539_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_16774_ clknet_leaf_117_wb_clk_i _02404_ _00470_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13986_ _07380_ _07468_ _03805_ vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__or3b_4
XTAP_TAPCELL_ROW_105_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09502__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15725_ net1265 vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__inv_2
X_12937_ net236 net2173 net470 vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13542__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10663__A2 _06125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15656_ net1248 vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_122_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12868_ net238 net2737 net478 vssd1 vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__mux2_1
XANTENNA__12666__B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14607_ net1239 vssd1 vssd1 vccd1 vccd1 _00237_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_174_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18375_ net1360 vssd1 vssd1 vccd1 vccd1 la_data_out[23] sky130_fd_sc_hd__buf_2
X_11819_ _07610_ _07615_ _07617_ vssd1 vssd1 vccd1 vccd1 _07631_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_174_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15587_ net1249 vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__inv_2
XANTENNA__08608__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12799_ net218 net2603 net487 vssd1 vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09678__D net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17326_ clknet_leaf_171_wb_clk_i _02956_ _01022_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14538_ net1121 vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__inv_2
XANTENNA__11612__B2 _07476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17257_ clknet_leaf_22_wb_clk_i _02887_ _00953_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14469_ net1185 vssd1 vssd1 vccd1 vccd1 _00099_ sky130_fd_sc_hd__inv_2
XANTENNA__10754__X _06753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16208_ net1216 vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17188_ clknet_leaf_181_wb_clk_i _02818_ _00884_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09033__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16139_ net1274 vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__inv_2
XANTENNA__08241__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10406__S net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08961_ _05017_ _05019_ _05021_ _05023_ vssd1 vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12621__S _03683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08892_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[17\]
+ net810 net736 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__a22o_1
XFILLER_0_166_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12628__A0 _03632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Left_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09513_ _05531_ net373 vssd1 vssd1 vccd1 vccd1 _05552_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_151_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11300__B1 _07129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13452__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15233__A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09444_ _05486_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[5\]
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_166_Right_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09375_ net375 _05419_ vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08326_ net948 net931 net925 vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__and3_1
XANTENNA__11603__B2 _07474_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09272__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08257_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[31\]
+ net701 net645 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[31\]
+ _04325_ vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__a221o_1
XANTENNA__09885__B _04533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08480__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout409_X net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08188_ _04237_ _04241_ _04231_ vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__a21oi_4
XANTENNA__09024__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout892_A _04279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_103_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10150_ net337 _06156_ _06163_ _06177_ vssd1 vssd1 vccd1 vccd1 _06178_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_37_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout680_X net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10590__A1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout778_X net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13627__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12531__S _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10081_ _04470_ _05998_ vssd1 vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10840__A team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12619__A0 _03657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13840_ net1456 net579 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[18\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_96_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13771_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[1\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[0\] team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[3\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[2\] vssd1
+ vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__or4_1
X_10983_ _06961_ _06962_ _06963_ net961 vssd1 vssd1 vccd1 vccd1 _06964_ sky130_fd_sc_hd__a211o_1
XANTENNA__08838__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13362__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15510_ net1167 vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12722_ _06737_ net1940 net499 vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16490_ clknet_leaf_182_wb_clk_i _02120_ _00186_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11390__B net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15441_ net1258 vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_133_Right_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12653_ net1610 _07350_ _03690_ vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_152_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11604_ net1601 net1010 net346 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03314_ sky130_fd_sc_hd__a22o_1
X_18160_ clknet_leaf_123_wb_clk_i _03463_ _01856_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15372_ net1078 vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__inv_2
X_12584_ net1677 _07791_ _03680_ vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_142_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09263__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17111_ clknet_leaf_145_wb_clk_i _02741_ _00807_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14323_ net375 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[7\]
+ _05442_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[6\] vssd1
+ vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__a22o_1
X_11535_ _07423_ _07428_ _07439_ _07445_ vssd1 vssd1 vccd1 vccd1 _07446_ sky130_fd_sc_hd__or4_2
X_18091_ clknet_leaf_67_wb_clk_i _03414_ _01787_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08471__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12706__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17042_ clknet_leaf_121_wb_clk_i _02672_ _00738_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input74_X net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14254_ _00023_ _00022_ _00038_ _00024_ vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__or4_1
Xwire375 _05397_ vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__buf_4
X_11466_ _07352_ _07371_ _07373_ _07376_ vssd1 vssd1 vccd1 vccd1 _07377_ sky130_fd_sc_hd__nand4_4
XANTENNA__09015__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13898__A2 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13205_ _06422_ net2928 net350 vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10417_ _05931_ _06056_ _06433_ net551 vssd1 vssd1 vccd1 vccd1 _06434_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_78_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14185_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[1\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__or2_1
X_11397_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[12\] _07327_
+ vssd1 vssd1 vccd1 vccd1 _07328_ sky130_fd_sc_hd__and2_1
XFILLER_0_150_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13136_ net230 net2121 net445 vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__mux2_1
X_10348_ _05980_ _05981_ vssd1 vssd1 vccd1 vccd1 _06368_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13537__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11846__A _07657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12441__S net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17944_ clknet_leaf_35_wb_clk_i _03283_ _01640_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10279_ net1021 _04677_ vssd1 vssd1 vccd1 vccd1 _06302_ sky130_fd_sc_hd__nand2_1
X_13067_ net242 net2422 net455 vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__mux2_1
X_12018_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[20\] team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[28\]
+ net993 _07518_ vssd1 vssd1 vccd1 vccd1 _07830_ sky130_fd_sc_hd__a31o_1
XANTENNA__10363__A2_N net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17875_ clknet_leaf_90_wb_clk_i _03218_ _01571_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10333__A1 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18350__1335 vssd1 vssd1 vccd1 vccd1 _18350__1335/HI net1335 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_124_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16826_ clknet_leaf_11_wb_clk_i _02456_ _00522_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_124_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16757_ clknet_leaf_24_wb_clk_i _02387_ _00453_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13969_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[7\] team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__nor2_1
XANTENNA__08829__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_181_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13272__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15708_ net1165 vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16688_ clknet_leaf_167_wb_clk_i _02318_ _00384_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15639_ net1245 vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09160_ _05211_ _05214_ _05210_ vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__and3b_1
XANTENNA__13586__A1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18358_ net1343 vssd1 vssd1 vccd1 vccd1 la_data_out[6] sky130_fd_sc_hd__buf_2
XFILLER_0_111_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09254__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08111_ net1028 net2451 vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__and2b_1
XFILLER_0_71_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17309_ clknet_leaf_109_wb_clk_i _02939_ _01005_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09091_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[12\]
+ net617 net614 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__a22o_1
XANTENNA__12616__S net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18289_ net1381 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
XANTENNA__08462__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08042_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[0\] vssd1
+ vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09006__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold901 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2315 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold912 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2326 sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2337 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold934 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold945 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold956 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net2392 sky130_fd_sc_hd__dlygate4sd3_1
Xhold989 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net2403 sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ _05350_ net365 vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__or2_1
XANTENNA__13447__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15228__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08944_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[16\]
+ net782 _05007_ net853 vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1013_A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08875_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[17\]
+ net711 net672 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[17\]
+ _04927_ vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_32_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout473_A _03706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout640_A net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13182__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout738_A _04421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09493__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09427_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[5\]
+ net689 net681 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[5\]
+ _05466_ vssd1 vssd1 vccd1 vccd1 _05470_ sky130_fd_sc_hd__a221o_1
XFILLER_0_109_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1170_X net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout905_A net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11037__C1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09358_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[7\]
+ net792 net775 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__a22o_1
XANTENNA__09245__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08309_ net1016 net943 net925 vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__and3_1
XFILLER_0_145_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12526__S net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09289_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[8\]
+ net693 net627 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[8\]
+ _05335_ vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__a221o_1
X_11320_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[112\] _07103_
+ _07105_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[8\] _07267_
+ vssd1 vssd1 vccd1 vccd1 _07279_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout895_X net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11251_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[51\] _07117_
+ _07121_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[83\] _07212_
+ vssd1 vssd1 vccd1 vccd1 _07213_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_56_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10202_ _06226_ _06227_ net527 vssd1 vssd1 vccd1 vccd1 _06228_ sky130_fd_sc_hd__mux2_1
X_11182_ _07141_ _07143_ _07145_ _07147_ vssd1 vssd1 vccd1 vccd1 _07148_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_128_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10133_ _06160_ vssd1 vssd1 vccd1 vccd1 _06161_ sky130_fd_sc_hd__inv_2
XANTENNA__13357__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15990_ net1130 vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_73_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input34_A gpio_in[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10064_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[14\] _06092_ vssd1
+ vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__and2_1
X_14941_ net1089 vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__inv_2
XANTENNA__10315__A1 _05634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17660_ clknet_leaf_77_wb_clk_i _03003_ _01356_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[98\]
+ sky130_fd_sc_hd__dfrtp_1
X_14872_ net1242 vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16611_ clknet_leaf_192_wb_clk_i _02241_ _00307_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13823_ net1543 net581 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[1\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_173_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17591_ clknet_leaf_73_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[28\]
+ _01287_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09469__C1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13092__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16542_ clknet_leaf_185_wb_clk_i _02172_ _00238_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13754_ _05212_ _06369_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[22\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__10618__A2 _06623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10966_ net1042 _06458_ vssd1 vssd1 vccd1 vccd1 _06950_ sky130_fd_sc_hd__nor2_1
XANTENNA__09484__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12705_ net255 net2285 net496 vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16473_ clknet_leaf_12_wb_clk_i _02103_ _00169_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11291__A2 _07105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08692__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13685_ net2887 net315 net386 vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__mux2_1
X_10897_ _06775_ _06776_ _06778_ _06885_ vssd1 vssd1 vccd1 vccd1 _06893_ sky130_fd_sc_hd__a211o_1
X_18212_ clknet_leaf_57_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.next_instr_wait
+ _01907_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.disable_pc
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15424_ net1113 vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__inv_2
X_12636_ _03605_ net1967 net201 vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09236__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18143_ clknet_leaf_126_wb_clk_i _03446_ _01839_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08444__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15355_ net1176 vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__inv_2
X_12567_ net2153 _07797_ _03678_ vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12436__S net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10745__A net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14306_ _04656_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[25\]
+ net379 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[24\] vssd1
+ vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__a22o_1
X_18074_ clknet_leaf_85_wb_clk_i _00015_ _01770_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11518_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read net1049
+ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[24\] vssd1 vssd1 vccd1
+ vccd1 _07429_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_124_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15286_ net1085 vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__inv_2
X_12498_ net1723 _07797_ _03673_ vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_117_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold208 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[30\] vssd1 vssd1
+ vccd1 vccd1 net1622 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_117_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold219 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[103\] vssd1 vssd1
+ vccd1 vccd1 net1633 sky130_fd_sc_hd__dlygate4sd3_1
X_17025_ clknet_leaf_151_wb_clk_i _02655_ _00721_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_14237_ _04023_ _04029_ vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__nor2_1
X_11449_ _07346_ _07359_ _07358_ vssd1 vssd1 vccd1 vccd1 _07360_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_169_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_169_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14168_ team_05_WB.instance_to_wrap.CPU_DAT_O\[17\] net504 net909 vssd1 vssd1 vccd1
+ vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[17\] sky130_fd_sc_hd__and3_1
XFILLER_0_21_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13267__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13119_ net303 net2575 net450 vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_84_Left_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12024__X _07836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14099_ _03950_ _03964_ vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__xnor2_1
X_17927_ clknet_leaf_43_wb_clk_i _03266_ _01623_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14887__A net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1270 net1271 vssd1 vssd1 vccd1 vccd1 net1270 sky130_fd_sc_hd__buf_4
XFILLER_0_56_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08660_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[23\]
+ net666 net649 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[23\]
+ _04722_ vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__a221o_1
Xfanout1281 net1312 vssd1 vssd1 vccd1 vccd1 net1281 sky130_fd_sc_hd__buf_2
X_17858_ clknet_leaf_91_wb_clk_i _03201_ _01554_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[40\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1292 net1294 vssd1 vssd1 vccd1 vccd1 net1292 sky130_fd_sc_hd__buf_4
XFILLER_0_89_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16809_ clknet_leaf_25_wb_clk_i _02439_ _00505_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_08591_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[25\]
+ net842 net791 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[25\]
+ _04666_ vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__a221o_1
X_17789_ clknet_leaf_101_wb_clk_i _03132_ _01485_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[99\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11515__S net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09475__A2 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_93_Left_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11282__A2 _07126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11019__C1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09212_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[10\]
+ net774 net752 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[10\]
+ _05263_ vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__a221o_1
XANTENNA__09227__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09143_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[11\]
+ net664 net640 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10242__B1 _04275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout319_A _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09074_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[13\]
+ net801 net760 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[13\]
+ _05126_ vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__a221o_1
XFILLER_0_114_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08025_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[31\] vssd1
+ vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1130_A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold720 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 net2145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold742 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2156 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1228_A net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold753 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2167 sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net2178 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout590_A _04368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold775 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net2189 sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2200 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13177__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout688_A net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold797 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 net2211 sky130_fd_sc_hd__dlygate4sd3_1
X_09976_ _05944_ _06004_ vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_51_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08927_ _04356_ _04991_ vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_51_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout855_A _04367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1420 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2834 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout476_X net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1431 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 net2845 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1442 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2856 sky130_fd_sc_hd__dlygate4sd3_1
X_08858_ _04923_ _04924_ vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__nor2_2
Xhold1453 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2867 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1464 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 net2878 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1475 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2889 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1486 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 net2900 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1497 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 net2911 sky130_fd_sc_hd__dlygate4sd3_1
X_08789_ net953 _04859_ _04346_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[19\]
+ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout643_X net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10820_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[12\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06817_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_49_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12470__A1 _07836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11273__A2 _07100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_98_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08674__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout810_X net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10751_ net332 _06613_ _06741_ _06749_ vssd1 vssd1 vccd1 vccd1 _06750_ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13640__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13470_ net226 net2309 net410 vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_27_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10682_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[5\] _06086_ vssd1
+ vssd1 vccd1 vccd1 _06685_ sky130_fd_sc_hd__or2_1
XANTENNA__09218__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_944 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12421_ _03632_ net1892 net215 vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08426__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10233__B1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15140_ net1229 vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__inv_2
X_12352_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[23\] team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[30\]
+ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[12\] net996 net545 vssd1
+ vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__a41o_1
XANTENNA__08035__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11303_ _07248_ _07249_ _07262_ vssd1 vssd1 vccd1 vccd1 _07263_ sky130_fd_sc_hd__or3_1
XFILLER_0_121_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15071_ net1178 vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_75_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12283_ _03568_ _03573_ _03576_ _03572_ vssd1 vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_75_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14022_ _03890_ _03891_ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11234_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[68\] _07118_
+ _07121_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[84\] _07196_
+ vssd1 vssd1 vccd1 vccd1 _07197_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_147_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10536__A1 _06049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_1_0_wb_clk_i_X clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13087__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11165_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[95\] _07096_
+ _07109_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[79\] vssd1 vssd1
+ vccd1 vccd1 _07131_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14278__A2 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10116_ _06142_ _06143_ vssd1 vssd1 vccd1 vccd1 _06144_ sky130_fd_sc_hd__nand2_1
X_11096_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[5\] _07062_
+ vssd1 vssd1 vccd1 vccd1 _07063_ sky130_fd_sc_hd__nor2_1
X_15973_ net1288 vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__inv_2
XANTENNA__09154__A1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[30\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17712_ clknet_leaf_93_wb_clk_i _03055_ _01408_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[86\]
+ sky130_fd_sc_hd__dfrtp_1
X_14924_ net1077 vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__inv_2
X_10047_ _06074_ _06075_ vssd1 vssd1 vccd1 vccd1 _06076_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_160_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold80 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[17\] vssd1 vssd1
+ vccd1 vccd1 net1494 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_160_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold91 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[19\]
+ vssd1 vssd1 vccd1 vccd1 net1505 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08901__A1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09153__X _05208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17643_ clknet_leaf_68_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[10\]
+ _01339_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_14855_ net1199 vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13806_ net2681 net971 net724 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[17\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_98_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17574_ clknet_leaf_113_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[11\]
+ _01270_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12020__A _07816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14786_ net1226 vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__inv_2
X_11998_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[17\] net995 _07724_
+ net548 vssd1 vssd1 vccd1 vccd1 _07810_ sky130_fd_sc_hd__a211o_1
XANTENNA__09457__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16525_ clknet_leaf_159_wb_clk_i _02155_ _00221_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13737_ net922 _06672_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[5\]
+ sky130_fd_sc_hd__nor2_1
X_10949_ _06795_ _06796_ _06873_ net1043 vssd1 vssd1 vccd1 vccd1 _06936_ sky130_fd_sc_hd__o31a_1
XANTENNA__12461__A1 _03604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08665__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13550__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16456_ clknet_leaf_197_wb_clk_i _02086_ _00152_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_119_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09209__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13668_ net2177 net229 net386 vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_119_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12674__B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15407_ net1138 vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12619_ _03657_ net1828 net202 vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__mux2_1
XANTENNA__13410__A0 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08417__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16387_ clknet_leaf_198_wb_clk_i _02017_ _00083_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13599_ net2060 net239 net395 vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09686__D net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18126_ clknet_leaf_48_wb_clk_i _00022_ _01822_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15338_ net1111 vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__inv_2
XANTENNA__09090__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10194__B _06219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18057_ net1037 _03395_ _01753_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[12\]
+ sky130_fd_sc_hd__dfrtp_4
X_15269_ net1203 vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__inv_2
XANTENNA__12690__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17008_ clknet_leaf_137_wb_clk_i _02638_ _00704_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout507 _07452_ vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09830_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[20\]
+ net841 net786 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__a22o_1
Xfanout518 net522 vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_158_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout529 net532 vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__clkbuf_4
X_09761_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[0\]
+ net663 _05771_ _05779_ _05788_ vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__a2111o_1
X_08712_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[22\]
+ net811 net783 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__a22o_1
X_09692_ _05721_ _05722_ _05723_ _05724_ vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__or4_1
XANTENNA__09696__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08643_ net379 _04716_ vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout269_A _06499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08574_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[25\]
+ net666 _04649_ net722 vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__a211o_1
XANTENNA__09448__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10369__B _05886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11255__A2 _07110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12452__A1 _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08656__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1080_A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout436_A _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08408__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout603_A net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09126_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[12\]
+ net786 _05181_ net853 vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__a211o_1
XFILLER_0_17_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09620__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09893__B _05921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09057_ _05109_ _05111_ _05113_ _05115_ vssd1 vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__or4_2
XANTENNA__12804__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_145_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_145_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold550 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net1964 sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[31\] vssd1 vssd1
+ vccd1 vccd1 net1975 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout593_X net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold572 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net1986 sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net1997 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1300_X net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold594 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2008 sky130_fd_sc_hd__dlygate4sd3_1
X_09959_ _05984_ _05987_ _05898_ vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout760_X net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13635__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12970_ net236 net2235 net466 vssd1 vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__mux2_1
Xhold1250 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2664 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09687__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1261 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 net2675 sky130_fd_sc_hd__dlygate4sd3_1
X_11921_ _07731_ _07732_ vssd1 vssd1 vccd1 vccd1 _07733_ sky130_fd_sc_hd__nand2_1
Xhold1272 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2686 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08895__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1283 net119 vssd1 vssd1 vccd1 vccd1 net2697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1294 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 net2708 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14640_ net1195 vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__inv_2
X_11852_ _07652_ _07662_ vssd1 vssd1 vccd1 vccd1 _07664_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_68_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[19\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[19\]
+ vssd1 vssd1 vccd1 vccd1 _06800_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12443__A1 _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11246__A2 _07097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08647__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14571_ net1073 vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__inv_2
X_11783_ _07573_ _07578_ _07591_ _07575_ vssd1 vssd1 vccd1 vccd1 _07595_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14319__X _04092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16310_ net1143 vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__inv_2
XANTENNA__13370__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13522_ net2782 net309 net404 vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17290_ clknet_leaf_3_wb_clk_i _02920_ _00986_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10734_ _06062_ _06733_ vssd1 vssd1 vccd1 vccd1 _06734_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16241_ net1144 vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_136_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13453_ net2456 net320 net414 vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__mux2_1
X_10665_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[6\] _06087_ vssd1
+ vssd1 vccd1 vccd1 _06669_ sky130_fd_sc_hd__xor2_1
XANTENNA__10295__A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08036__Y _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_149_Left_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12404_ _07840_ _07850_ _07851_ vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__and3_4
X_16172_ net1152 vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__inv_2
X_13384_ net1968 net300 net422 vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__mux2_1
XANTENNA__09072__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10596_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[10\] net905 net896
+ _06603_ vssd1 vssd1 vccd1 vccd1 _06604_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_51_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10757__A1 _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15123_ net1212 vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__inv_2
X_12335_ _03627_ _03628_ _03629_ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_11_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12714__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15054_ net1187 vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12266_ _03555_ _03556_ vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__nand2b_1
X_14005_ _03850_ _03875_ vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_142_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11217_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[5\] _07100_ _07104_
+ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[117\] _07180_ vssd1
+ vssd1 vccd1 vccd1 _07181_ sky130_fd_sc_hd__a221o_1
X_12197_ _08004_ _08006_ _07999_ vssd1 vssd1 vccd1 vccd1 _08009_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08212__B net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_162_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__clkbuf_4
X_11148_ _07072_ _07088_ vssd1 vssd1 vccd1 vccd1 _07114_ sky130_fd_sc_hd__or2_4
XPHY_EDGE_ROW_158_Left_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13545__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15326__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11079_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[0\] _07032_
+ _07043_ _07045_ vssd1 vssd1 vccd1 vccd1 _07046_ sky130_fd_sc_hd__a211o_1
X_15956_ net1307 vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__inv_2
XANTENNA__12669__B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14907_ net1176 vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__inv_2
X_15887_ net1302 vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08350__A2 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17626_ clknet_leaf_62_wb_clk_i _02997_ _01322_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10693__B1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14838_ net1101 vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11237__A2 _07115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17557_ clknet_leaf_59_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[28\]
+ _01253_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_14769_ net1189 vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__inv_2
XANTENNA__08638__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08102__A2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[10\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13280__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16508_ clknet_leaf_156_wb_clk_i _02138_ _00204_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_17488_ clknet_leaf_37_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[23\]
+ _01184_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_08290_ _04236_ _04240_ _04150_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[20\]
+ _04230_ vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_129_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09850__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[20\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_167_Left_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16439_ clknet_leaf_145_wb_clk_i _02069_ _00135_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17984__Q net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18109_ clknet_leaf_55_wb_clk_i _03432_ _01805_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12624__S net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout304 _06655_ vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout315 net316 vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__buf_2
XANTENNA__08574__C1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout326 net327 vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__clkbuf_2
Xfanout337 _06050_ vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__clkbuf_4
X_09813_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[20\]
+ net664 net644 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__a22o_1
Xfanout348 _06063_ vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout359 _07296_ vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__buf_2
XANTENNA_fanout386_A net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13455__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09744_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[0\]
+ net880 net861 net859 vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__and4_1
XANTENNA__09669__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09675_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[1\]
+ net876 net864 net862 vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__and4_1
XANTENNA__08341__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10684__B1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08626_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[24\]
+ net812 net746 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11228__A2 _07103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08557_ _04613_ _04632_ vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__or2_1
XANTENNA__08629__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout720_A _04285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout341_X net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout439_X net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout818_A net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13190__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08488_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[27\]
+ net666 net661 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__a22o_1
XANTENNA__09841__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18282__A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout606_X net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10450_ net892 _06464_ vssd1 vssd1 vccd1 vccd1 _06465_ sky130_fd_sc_hd__nor2_1
XANTENNA__09054__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11498__X _07409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09109_ _04158_ _04353_ vssd1 vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11939__A team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12534__S net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10381_ _06394_ _06399_ net538 vssd1 vssd1 vccd1 vccd1 _06400_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08801__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12120_ _07927_ _07929_ vssd1 vssd1 vccd1 vccd1 _07932_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08313__A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12051_ _07363_ _07860_ _07862_ vssd1 vssd1 vccd1 vccd1 _07863_ sky130_fd_sc_hd__a21oi_4
Xhold380 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[118\] vssd1 vssd1
+ vccd1 vccd1 net1794 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold391 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[83\] vssd1 vssd1
+ vccd1 vccd1 net1805 sky130_fd_sc_hd__dlygate4sd3_1
X_11002_ _06858_ _06978_ vssd1 vssd1 vccd1 vccd1 _06979_ sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_leaf_59_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_99_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14321__Y _04094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout860 net861 vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__buf_2
XANTENNA__13365__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15810_ net1298 vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__inv_2
XANTENNA__08580__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout871 net873 vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__buf_2
X_16790_ clknet_leaf_138_wb_clk_i _02420_ _00486_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout882 _04282_ vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__clkbuf_2
Xfanout893 net894 vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__buf_2
X_15741_ net1269 vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__inv_2
X_12953_ net294 net2421 net470 vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__mux2_1
XANTENNA__08868__B1 _04314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1080 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2494 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_172_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1091 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 net2505 sky130_fd_sc_hd__dlygate4sd3_1
X_11904_ _07681_ _07715_ net343 vssd1 vssd1 vccd1 vccd1 _07716_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_107_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15672_ net1259 vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_42_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_66_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ net300 net2073 net477 vssd1 vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__mux2_1
X_17411_ clknet_leaf_65_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[11\]
+ _01107_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_14623_ net1184 vssd1 vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__inv_2
XANTENNA__11219__A2 _07113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18391_ net1370 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__buf_2
X_11835_ _07590_ _07646_ _07639_ vssd1 vssd1 vccd1 vccd1 _07647_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_157_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12709__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17342_ clknet_leaf_40_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[6\]
+ _01038_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_14554_ net1052 vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__inv_2
X_11766_ _07548_ _07560_ vssd1 vssd1 vccd1 vccd1 _07578_ sky130_fd_sc_hd__or2_1
XANTENNA__09293__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10978__A1 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09832__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10737__B _06736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ net2466 net253 net404 vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__mux2_1
X_10717_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[3\] team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06718_ sky130_fd_sc_hd__or2_1
X_17273_ clknet_leaf_12_wb_clk_i _02903_ _00969_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14485_ net1079 vssd1 vssd1 vccd1 vccd1 _00115_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11697_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[19\] team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[21\]
+ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[23\] team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[30\]
+ net993 vssd1 vssd1 vccd1 vccd1 _07509_ sky130_fd_sc_hd__o41a_1
XANTENNA__08207__B net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16224_ net1228 vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__inv_2
X_13436_ net2715 net232 net415 vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10648_ _06088_ _06652_ vssd1 vssd1 vccd1 vccd1 _06653_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_24_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08399__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14325__A2_N _05768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16155_ net1253 vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_98_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12444__S net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13367_ net2788 net243 net422 vssd1 vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__mux2_1
X_10579_ _06585_ _06587_ _04264_ vssd1 vssd1 vccd1 vccd1 _06588_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_24_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15106_ net1226 vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12318_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[18\] net996 _03586_
+ net545 vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__a211o_1
XFILLER_0_11_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16086_ net1308 vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__inv_2
X_13298_ net2589 net190 net430 vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15037_ net1088 vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__inv_2
X_12249_ _08019_ _03543_ vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__or2_1
XANTENNA__14341__B2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13275__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08571__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16988_ clknet_leaf_157_wb_clk_i _02618_ _00684_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_147_Right_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15939_ net1304 vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__inv_2
XANTENNA__08859__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08323__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10666__B1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09460_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[5\]
+ _04366_ net828 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[5\]
+ net856 vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__a221o_1
XANTENNA__09989__A _05208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08411_ _04490_ vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__inv_2
X_17609_ clknet_leaf_66_wb_clk_i _02980_ _01305_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_09391_ _05430_ _05432_ _05433_ _05435_ vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__or4_2
XANTENNA__12619__S net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10418__B1 _06355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08342_ _04405_ _04410_ _04416_ _04423_ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__or4_1
XANTENNA__09284__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09823__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08273_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[16\] team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[15\]
+ _04355_ vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_15_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09036__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12040__C1 _07840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout301_A _06621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1043_A net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1210_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11697__A2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[21\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout670_A net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13185__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08562__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout768_A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout389_X net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout189 net192 vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09727_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[0\]
+ net745 _05744_ _05745_ _05755_ vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__a2111oi_1
XTAP_TAPCELL_ROW_87_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout935_A net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout556_X net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09658_ _05688_ _05689_ _05690_ _05691_ vssd1 vssd1 vccd1 vccd1 _05692_ sky130_fd_sc_hd__or4_1
XFILLER_0_167_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08609_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[24\]
+ net697 net642 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[24\]
+ _04683_ vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__a221o_1
XANTENNA__12529__S net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09589_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[2\]
+ net846 _05600_ _05606_ _05617_ vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10838__A team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11620_ net2934 net1010 net345 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__a22o_1
XANTENNA__09275__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09814__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08308__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_132_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_108_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11551_ _07398_ _07459_ _07460_ _07461_ vssd1 vssd1 vccd1 vccd1 _07462_ sky130_fd_sc_hd__nand4_1
XANTENNA__12475__D _03659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10502_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[15\] _06093_ vssd1
+ vssd1 vccd1 vccd1 _06515_ sky130_fd_sc_hd__xnor2_1
X_14270_ _04043_ _04048_ vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire535 _05234_ vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__buf_4
XANTENNA__09027__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11482_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[25\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[25\]
+ net1034 vssd1 vssd1 vccd1 vccd1 _07393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_160_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_160_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_45_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13221_ net2024 net353 vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_150_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10433_ _06448_ vssd1 vssd1 vccd1 vccd1 _06449_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_150_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12582__A0 _03651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input64_A wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13152_ net302 net2704 net445 vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__mux2_1
X_10364_ net895 _06382_ _06383_ _05259_ vssd1 vssd1 vccd1 vccd1 _06384_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_103_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12103_ _07902_ _07909_ _07912_ _07907_ vssd1 vssd1 vccd1 vccd1 _07915_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_130_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14323__A1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13083_ net288 net2557 net452 vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__mux2_1
XANTENNA__14323__B2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17960_ clknet_leaf_107_wb_clk_i _03299_ _01656_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__dfrtp_1
X_10295_ net383 _06317_ vssd1 vssd1 vccd1 vccd1 _06318_ sky130_fd_sc_hd__and2_1
X_12034_ _07365_ net919 _07352_ vssd1 vssd1 vccd1 vccd1 _07846_ sky130_fd_sc_hd__o21a_1
X_16911_ clknet_leaf_141_wb_clk_i _02541_ _00607_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_17891_ clknet_leaf_76_wb_clk_i _03234_ _01587_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13095__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08553__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16842_ clknet_leaf_194_wb_clk_i _02472_ _00538_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_109_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout690 _04299_ vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__buf_4
X_13985_ _03855_ _03856_ vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__nor2_1
X_16773_ clknet_leaf_18_wb_clk_i _02403_ _00469_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_171_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_73_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15724_ net1299 vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__inv_2
X_12936_ net239 net2594 net470 vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15655_ net1248 vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__inv_2
X_12867_ net243 net2143 net478 vssd1 vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_122_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14606_ net1189 vssd1 vssd1 vccd1 vccd1 _00236_ sky130_fd_sc_hd__inv_2
X_11818_ _07615_ _07617_ _07610_ vssd1 vssd1 vccd1 vccd1 _07630_ sky130_fd_sc_hd__a21boi_2
X_18374_ net1359 vssd1 vssd1 vccd1 vccd1 la_data_out[22] sky130_fd_sc_hd__buf_2
X_15586_ net1250 vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__inv_2
XANTENNA__09266__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12798_ net189 net2388 net485 vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_174_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_174_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17325_ clknet_leaf_162_wb_clk_i _02955_ _01021_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[21\]
+ sky130_fd_sc_hd__dfrtp_2
X_14537_ net1221 vssd1 vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__inv_2
X_11749_ _07560_ vssd1 vssd1 vccd1 vccd1 _07561_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17256_ clknet_leaf_203_wb_clk_i _02886_ _00952_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_14468_ net1230 vssd1 vssd1 vccd1 vccd1 _00098_ sky130_fd_sc_hd__inv_2
XANTENNA__12682__B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13419_ net2055 net304 net418 vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__mux2_1
X_16207_ net1184 vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__inv_2
X_17187_ clknet_leaf_191_wb_clk_i _02817_ _00883_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_14399_ net1533 vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12573__A0 _03650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16138_ net1274 vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08792__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16069_ net1260 vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__inv_2
X_08960_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[15\]
+ net648 net598 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[15\]
+ _05022_ vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__a221o_1
XANTENNA__12902__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08891_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[17\]
+ net841 net821 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[17\]
+ _04956_ vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__a221o_1
XANTENNA__08544__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09512_ net373 _05531_ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_91_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09443_ _04246_ _04349_ _05484_ _05485_ vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_82_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10658__A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09374_ net573 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[7\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[7\] vssd1 vssd1 vccd1
+ vccd1 _05419_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08325_ _04270_ net1017 net951 net938 vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11603__A2 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1160_A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1258_A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08256_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[31\]
+ net684 net613 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[31\]
+ _04324_ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09009__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08187_ _04237_ _04241_ _04231_ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__a21o_2
XANTENNA__12564__A0 _03664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_104_Left_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout885_A _04281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12812__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1213_X net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10080_ _04470_ _05919_ vssd1 vssd1 vccd1 vccd1 _06108_ sky130_fd_sc_hd__xnor2_4
XTAP_TAPCELL_ROW_89_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout673_X net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14312__B _04084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12113__A _07914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout840_X net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout938_X net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Left_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13643__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13770_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[5\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[4\] team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[7\]
+ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[6\] vssd1
+ vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__or4_1
X_10982_ net1043 _06515_ vssd1 vssd1 vccd1 vccd1 _06963_ sky130_fd_sc_hd__nor2_1
XANTENNA__09496__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12721_ net312 net2135 net496 vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10568__A _06049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15440_ net1253 vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12652_ _03687_ _03689_ vssd1 vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_100_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09248__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11603_ net1719 net1010 _07472_ _07474_ vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__a22o_1
X_15371_ net1077 vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_152_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12583_ net1715 _07789_ _03680_ vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__mux2_1
X_17110_ clknet_leaf_140_wb_clk_i _02740_ _00806_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14322_ _04990_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__nor2_1
X_11534_ _07357_ _07360_ _07441_ _07444_ vssd1 vssd1 vccd1 vccd1 _07445_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_151_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18090_ clknet_leaf_79_wb_clk_i _03413_ _01786_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_122_Left_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17041_ clknet_leaf_172_wb_clk_i _02671_ _00737_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14253_ _00021_ team_05_WB.instance_to_wrap.total_design.keypad0.counter\[1\] _04036_
+ _04037_ vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__or4_1
X_11465_ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[5\] _07375_ net1002
+ vssd1 vssd1 vccd1 vccd1 _07376_ sky130_fd_sc_hd__mux2_2
XFILLER_0_80_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12555__A0 _03610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwire376 _04900_ vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__buf_4
XFILLER_0_123_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13204_ _06404_ net2713 net350 vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10416_ net1018 _04881_ _04879_ vssd1 vssd1 vccd1 vccd1 _06433_ sky130_fd_sc_hd__o21a_1
X_14184_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[0\] net729
+ vssd1 vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__and2b_1
XFILLER_0_151_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11396_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[11\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[10\]
+ _07326_ vssd1 vssd1 vccd1 vccd1 _07327_ sky130_fd_sc_hd__and3_1
XANTENNA__09420__B1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08774__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13135_ net235 net2328 net446 vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10347_ net2211 net230 net541 vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__mux2_1
XANTENNA__12722__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13066_ net224 net2555 net454 vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__mux2_1
X_17943_ clknet_leaf_33_wb_clk_i _03282_ _01639_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10278_ _06003_ _06300_ vssd1 vssd1 vccd1 vccd1 _06301_ sky130_fd_sc_hd__nor2_1
X_12017_ _07515_ _07530_ _07828_ vssd1 vssd1 vccd1 vccd1 _07829_ sky130_fd_sc_hd__and3_1
XANTENNA__08526__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17874_ clknet_leaf_92_wb_clk_i _03217_ _01570_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08220__B net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16825_ clknet_leaf_10_wb_clk_i _02455_ _00521_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_124_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13553__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12310__X _03605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09487__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16756_ clknet_leaf_119_wb_clk_i _02386_ _00452_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13968_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[7\] team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__and2_1
XANTENNA__12677__B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15707_ net1166 vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__inv_2
XANTENNA__11294__B1 _07124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12919_ net303 net2277 net474 vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__mux2_1
X_13899_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[21\]
+ net558 net574 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[21\]
+ net985 vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__a221o_1
X_16687_ clknet_leaf_134_wb_clk_i _02317_ _00383_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09239__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15638_ net1281 vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18357_ net1342 vssd1 vssd1 vccd1 vccd1 la_data_out[5] sky130_fd_sc_hd__buf_2
XFILLER_0_28_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15569_ net1246 vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__inv_2
X_08110_ net1029 net1022 net975 _04204_ vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11597__B2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[27\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17308_ clknet_leaf_154_wb_clk_i _02938_ _01004_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09090_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[12\]
+ net676 net668 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18288_ net1380 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
XANTENNA__08235__X _04318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08041_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[3\] vssd1
+ vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17239_ clknet_leaf_144_wb_clk_i _02869_ _00935_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12546__A0 _03661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold902 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2316 sky130_fd_sc_hd__dlygate4sd3_1
Xhold913 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net2327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold924 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2338 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09411__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_83 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold935 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold946 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2382 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12632__S net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09992_ net349 net365 vssd1 vssd1 vccd1 vccd1 _06021_ sky130_fd_sc_hd__nand2_1
Xhold979 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 net2393 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08943_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[16\]
+ net802 net748 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__a22o_1
XANTENNA__08411__A _04490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09175__C1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout299_A _06621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08874_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[17\]
+ net594 _04940_ net720 vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_32_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11521__A1 _07346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10324__A2 _06345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09190__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout466_A _03710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13463__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15244__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09478__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10088__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout633_A _04313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09426_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[5\]
+ net623 net616 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09357_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[7\]
+ net842 net769 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout421_X net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12807__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout800_A net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1163_X net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11588__A1 _07354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11588__B2 net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08308_ net1015 net949 net925 vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__and3_1
XFILLER_0_62_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09288_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[8\]
+ net681 net631 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[8\]
+ _05336_ vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__a221o_1
XFILLER_0_118_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08239_ net884 net874 net861 vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__and3_1
XFILLER_0_166_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12537__A0 _07816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08305__B net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11250_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[27\] _07119_
+ _07120_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[35\] vssd1 vssd1
+ vccd1 vccd1 _07212_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09402__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout790_X net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout888_X net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13638__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10201_ _06128_ _06138_ net518 vssd1 vssd1 vccd1 vccd1 _06227_ sky130_fd_sc_hd__mux2_1
XANTENNA__08756__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11181_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[119\] _07104_
+ _07106_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[23\] _07146_
+ vssd1 vssd1 vccd1 vccd1 _07147_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_128_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10132_ net524 _06159_ vssd1 vssd1 vccd1 vccd1 _06160_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08508__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10063_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[13\] team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[12\]
+ _06091_ vssd1 vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__and3_1
X_14940_ net1095 vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_145_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09704__X team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input27_A DAT_I[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14871_ net1099 vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_1030 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13373__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16610_ clknet_leaf_4_wb_clk_i _02240_ _00306_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13822_ net1474 net578 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_write_data\[0\]
+ sky130_fd_sc_hd__and2_1
X_17590_ clknet_leaf_113_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[27\]
+ _01286_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11276__B1 _07118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13753_ net921 _06387_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[21\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16541_ clknet_leaf_131_wb_clk_i _02171_ _00237_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10965_ _06802_ _06803_ _06805_ _06868_ vssd1 vssd1 vccd1 vccd1 _06949_ sky130_fd_sc_hd__a211o_1
XFILLER_0_35_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12704_ net253 net2572 net496 vssd1 vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13684_ net1998 net317 net385 vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__mux2_1
X_16472_ clknet_leaf_27_wb_clk_i _02102_ _00168_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10896_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[31\] net565 _06891_
+ _06892_ vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18211_ clknet_leaf_50_wb_clk_i net1416 _01906_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_fetch
+ sky130_fd_sc_hd__dfrtp_4
X_12635_ net1669 _07797_ _03682_ vssd1 vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__mux2_1
X_15423_ net1114 vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__inv_2
XANTENNA__12717__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_130_Left_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15354_ net1056 vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__inv_2
X_18142_ clknet_leaf_151_wb_clk_i _03445_ _01838_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12566_ net1773 _07798_ _03678_ vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10745__B _06743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11517_ _07425_ _07427_ net920 vssd1 vssd1 vccd1 vccd1 _07428_ sky130_fd_sc_hd__o21a_1
X_14305_ _04077_ vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__inv_2
X_18073_ clknet_leaf_85_wb_clk_i _00014_ _01769_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_15285_ net1060 vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__inv_2
XANTENNA__12528__A0 _03663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12497_ net1703 _07798_ _03673_ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14236_ team_05_WB.instance_to_wrap.total_design.keypad0.counter\[10\] _04022_ net2474
+ vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__a21oi_1
Xhold209 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[41\] vssd1 vssd1
+ vccd1 vccd1 net1623 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17024_ clknet_leaf_129_wb_clk_i _02654_ _00720_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11448_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[29\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[29\]
+ net1033 vssd1 vssd1 vccd1 vccd1 _07359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_169_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11200__B1 _07116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08747__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13548__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12452__S net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14167_ net2971 net502 net908 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[16\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__15329__A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11379_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[1\] _07052_
+ net731 vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__mux2_1
XANTENNA__10554__A2 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13118_ net295 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[8\]
+ net451 vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__mux2_1
X_14098_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[15\] net978 team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[13\]
+ _04160_ vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__o31a_1
X_17926_ clknet_leaf_43_wb_clk_i _03265_ _01622_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13049_ net292 net2707 net456 vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1260 net1261 vssd1 vssd1 vccd1 vccd1 net1260 sky130_fd_sc_hd__clkbuf_4
Xfanout1271 net1279 vssd1 vssd1 vccd1 vccd1 net1271 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09172__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17857_ clknet_leaf_100_wb_clk_i _03200_ _01553_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[39\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1282 net1283 vssd1 vssd1 vccd1 vccd1 net1282 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_1_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1293 net1294 vssd1 vssd1 vccd1 vccd1 net1293 sky130_fd_sc_hd__buf_4
XANTENNA__08380__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13283__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16808_ clknet_leaf_1_wb_clk_i _02438_ _00504_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12040__X _07852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08590_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[25\]
+ net811 net761 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__a22o_1
X_17788_ clknet_leaf_77_wb_clk_i _03131_ _01484_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[98\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11267__B1 _07109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16739_ clknet_leaf_198_wb_clk_i _02369_ _00435_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09997__A _05078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09211_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[10\]
+ net821 net802 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__a22o_1
X_18409_ net913 vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12627__S net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09142_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[11\]
+ net648 net632 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[11\]
+ _05196_ vssd1 vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__a221o_1
XANTENNA__13964__C1 _07451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08986__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09073_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[13\]
+ net836 net826 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[13\]
+ _05127_ vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__a221o_1
XFILLER_0_170_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout214_A net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold710 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold721 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2135 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold732 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 net2146 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13192__A0 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08738__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13458__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold743 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 net2157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold754 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net2168 sky130_fd_sc_hd__dlygate4sd3_1
Xhold765 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold776 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2190 sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net2201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold798 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2212 sky130_fd_sc_hd__dlygate4sd3_1
X_09975_ _05731_ net362 vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__or2_1
XANTENNA__09148__C1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08926_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[15\] _04355_
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[16\] vssd1 vssd1
+ vccd1 vccd1 _04991_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_51_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1410 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2824 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09163__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1421 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2835 sky130_fd_sc_hd__dlygate4sd3_1
X_08857_ net376 _04921_ vssd1 vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__and2_1
Xhold1432 net132 vssd1 vssd1 vccd1 vccd1 net2846 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout750_A net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1443 team_05_WB.instance_to_wrap.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 net2857
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1454 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2868 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1465 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2879 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08371__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout848_A _04373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout469_X net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08910__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1476 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 net2890 sky130_fd_sc_hd__dlygate4sd3_1
X_08788_ _04152_ _04358_ vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__xnor2_1
Xhold1487 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2901 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_140_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1498 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net2912 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11258__B1 _07128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1280_X net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout636_X net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15702__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10750_ _06747_ _06748_ _06745_ vssd1 vssd1 vccd1 vccd1 _06749_ sky130_fd_sc_hd__a21oi_1
X_09409_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[6\]
+ net806 net746 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[6\]
+ _05452_ vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__a221o_1
XFILLER_0_165_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12537__S _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10681_ _06675_ _06682_ _06683_ net537 vssd1 vssd1 vccd1 vccd1 _06684_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout803_X net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10846__A team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12420_ _03612_ net1856 net214 vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10233__A1 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12351_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[23\] net1000 net546
+ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__a21o_2
XANTENNA__08977__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_67_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_63_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11302_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[41\] _07091_
+ _07092_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[1\] _07261_
+ vssd1 vssd1 vccd1 vccd1 _07262_ sky130_fd_sc_hd__a221o_1
X_15070_ net1063 vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12282_ _07986_ _03575_ vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14021_ _03887_ _03889_ vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__and2_1
XANTENNA__13368__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11233_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[76\] _07116_
+ _07119_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[28\] vssd1 vssd1
+ vccd1 vccd1 _07196_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_858 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08729__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11164_ _07068_ _07071_ _07079_ vssd1 vssd1 vccd1 vccd1 _07130_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_112_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14988__A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10115_ _04944_ net367 vssd1 vssd1 vccd1 vccd1 _06143_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_164_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11095_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[3\] _07061_
+ _07034_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[4\] vssd1
+ vssd1 vccd1 vccd1 _07062_ sky130_fd_sc_hd__o2bb2a_1
X_15972_ net1293 vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__inv_2
X_17711_ clknet_leaf_86_wb_clk_i _03054_ _01407_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[85\]
+ sky130_fd_sc_hd__dfrtp_1
X_14923_ net1070 vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__inv_2
X_10046_ _04613_ net367 vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__nor2_1
XANTENNA__08898__D1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold70 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[30\]
+ vssd1 vssd1 vccd1 vccd1 net1484 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08362__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold81 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[28\]
+ vssd1 vssd1 vccd1 vccd1 net1495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[13\]
+ vssd1 vssd1 vccd1 vccd1 net1506 sky130_fd_sc_hd__dlygate4sd3_1
X_17642_ clknet_leaf_68_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[9\]
+ _01338_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08901__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[17\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14854_ net1247 vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__inv_2
XANTENNA__11249__B1 _07169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13805_ net1593 net970 net723 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[16\]
+ sky130_fd_sc_hd__and3_1
X_17573_ clknet_leaf_113_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[10\]
+ _01269_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11997_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[18\] net995 _07722_
+ net548 vssd1 vssd1 vccd1 vccd1 _07809_ sky130_fd_sc_hd__a211o_1
X_14785_ net1235 vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12795__X _03703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16524_ clknet_leaf_0_wb_clk_i _02154_ _00220_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13736_ net923 _06691_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[4\]
+ sky130_fd_sc_hd__nor2_1
X_10948_ _06795_ _06796_ _06873_ vssd1 vssd1 vccd1 vccd1 _06935_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10472__A1 _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16455_ clknet_leaf_200_wb_clk_i _02085_ _00151_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10879_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[22\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[22\]
+ _06875_ vssd1 vssd1 vccd1 vccd1 _06876_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12447__S net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13667_ net2680 net233 net385 vssd1 vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_119_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15406_ net1133 vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__inv_2
X_12618_ net1768 _07791_ _03682_ vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16386_ clknet_leaf_5_wb_clk_i _02016_ _00082_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13598_ net1972 net243 net395 vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18125_ clknet_leaf_48_wb_clk_i _00039_ _01821_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08968__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12549_ net1858 _07789_ _03678_ vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15337_ net1225 vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18056_ net1037 _03394_ _01752_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_1 _06518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15268_ net1237 vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__inv_2
XANTENNA__13278__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17007_ clknet_leaf_141_wb_clk_i _02637_ _00703_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_14219_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[13\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[14\]
+ _04013_ vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__nand3_1
XANTENNA__15059__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15199_ net1182 vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__inv_2
XANTENNA__09393__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout508 net509 vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__buf_2
XFILLER_0_67_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout519 net522 vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__clkbuf_2
X_09760_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[0\]
+ net620 _05774_ _05775_ _05778_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12910__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08711_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[22\]
+ net820 _04783_ vssd1 vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__a21o_1
X_17909_ clknet_leaf_103_wb_clk_i _03252_ _01605_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09145__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09691_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[1\]
+ net690 _05703_ _05704_ _05718_ vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08353__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11526__S net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1090 net1094 vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__clkbuf_4
X_08642_ net570 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[24\]
+ _04362_ vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__o21a_1
XFILLER_0_83_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08573_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[25\]
+ net654 net609 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15522__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10463__A1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout331_A _06705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17510__Q team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout429_A net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10385__B _06403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09125_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[12\]
+ net833 net793 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08959__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout217_X net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1240_A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10766__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09056_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[13\]
+ net607 net598 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[13\]
+ _05114_ vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__a221o_1
XFILLER_0_170_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08158__A_N team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13188__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout798_A net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold540 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net1954 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold551 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[14\] vssd1
+ vssd1 vccd1 vccd1 net1965 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10518__A2 _06525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold562 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 net1976 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09384__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold573 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 net1987 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_49_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_130_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold584 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net1998 sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 net100 vssd1 vssd1 vccd1 vccd1 net2009 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11191__A2 _07124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08592__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08302__C net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12820__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09958_ _05929_ _05986_ _05985_ vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_185_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_185_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_142_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09136__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08909_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[16\]
+ net691 net683 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[16\]
+ _04972_ vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout753_X net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09889_ _04554_ _05917_ vssd1 vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__nand2_2
XANTENNA__14320__B team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[15\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_114_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_114_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold1240 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1251 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[9\] vssd1 vssd1
+ vccd1 vccd1 net2665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1262 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2676 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11920_ _07695_ _07697_ vssd1 vssd1 vccd1 vccd1 _07732_ sky130_fd_sc_hd__nand2b_1
Xhold1273 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net2687 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1284 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 net2698 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1295 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net2709 sky130_fd_sc_hd__dlygate4sd3_1
X_11851_ _07652_ _07662_ vssd1 vssd1 vccd1 vccd1 _07663_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout920_X net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13651__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ _06797_ _06798_ vssd1 vssd1 vccd1 vccd1 _06799_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14570_ net1121 vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__inv_2
X_11782_ _07585_ _07588_ _07591_ _07592_ _07582_ vssd1 vssd1 vccd1 vccd1 _07594_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_28_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09844__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13521_ net2690 net329 net406 vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__mux2_1
X_10733_ _06596_ _06726_ net370 vssd1 vssd1 vccd1 vccd1 _06733_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16240_ net1135 vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13452_ net1957 net304 net414 vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__mux2_1
X_10664_ _06659_ _06660_ _06667_ net537 vssd1 vssd1 vccd1 vccd1 _06668_ sky130_fd_sc_hd__a31o_1
XFILLER_0_119_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10295__B _06317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12403_ net1695 _03623_ net217 vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16171_ net1143 vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__inv_2
X_13383_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[10\]
+ net286 net420 vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_88_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10595_ _06090_ _06602_ vssd1 vssd1 vccd1 vccd1 _06603_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16344__RESET_B _00040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12334_ net354 _03598_ _03626_ _03616_ _07512_ vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_114_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15122_ net1232 vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13098__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15053_ net1081 vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__inv_2
X_12265_ _03559_ vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14004_ _03872_ _03873_ vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__xor2_1
XFILLER_0_120_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11216_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[93\] _07108_
+ _07129_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[61\] vssd1 vssd1
+ vccd1 vccd1 _07180_ sky130_fd_sc_hd__a22o_1
X_12196_ _08004_ _08006_ vssd1 vssd1 vccd1 vccd1 _08008_ sky130_fd_sc_hd__nand2_1
XANTENNA__08583__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__clkbuf_4
XANTENNA__08212__C net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 ADR_O[26] sky130_fd_sc_hd__clkbuf_4
X_11147_ _07074_ _07112_ vssd1 vssd1 vccd1 vccd1 _07113_ sky130_fd_sc_hd__nor2_4
XANTENNA__12730__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09127__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11078_ _04164_ _07044_ vssd1 vssd1 vccd1 vccd1 _07045_ sky130_fd_sc_hd__and2_1
X_15955_ net1303 vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__inv_2
X_14906_ net1058 vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__inv_2
X_10029_ net381 net364 vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__nor2_1
X_15886_ net1272 vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__inv_2
X_17625_ clknet_leaf_59_wb_clk_i _02996_ _01321_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_14837_ net1079 vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__inv_2
XANTENNA__13561__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15342__A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17556_ clknet_leaf_65_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[27\]
+ _01252_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09835__B1 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14768_ net1183 vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12685__B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16507_ clknet_leaf_191_wb_clk_i _02137_ _00203_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13719_ net905 _06424_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[19\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_74_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17487_ clknet_leaf_37_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[22\]
+ _01183_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_14699_ net1070 vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16438_ clknet_leaf_142_wb_clk_i _02068_ _00134_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12905__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16369_ clknet_leaf_122_wb_clk_i _01999_ _00065_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_18108_ clknet_leaf_55_wb_clk_i _03431_ _01804_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[25\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_143_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18039_ clknet_leaf_96_wb_clk_i _03377_ _01735_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_23_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13698__A1 team_05_WB.instance_to_wrap.wishbone.curr_state\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout305 net308 vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11173__A2 _07125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout316 _06688_ vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12370__A1 _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09812_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[20\]
+ net691 net621 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__a22o_1
Xfanout327 _06753_ vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__buf_2
XANTENNA__12640__S _03682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout338 _06050_ vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10381__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09118__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09743_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[0\]
+ net886 net868 net863 vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__and4_1
XFILLER_0_20_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09674_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[1\]
+ net876 net874 net862 vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__and4_1
XFILLER_0_55_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10684__A1 _04173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08625_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[24\]
+ net758 net742 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1190_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout546_A _07467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13471__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08556_ net570 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[26\]
+ _04362_ vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_46_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13622__A1 _06737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10667__Y _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09826__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10436__A1 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_122_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08487_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[27\]
+ net701 net608 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[27\]
+ _04564_ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__a221o_1
XFILLER_0_64_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout334_X net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout713_A _04288_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1243_X net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12815__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09108_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[12\]
+ net715 _05160_ _05164_ vssd1 vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__o22ai_4
X_10380_ net555 _06390_ _06398_ net348 vssd1 vssd1 vccd1 vccd1 _06399_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_131_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_14_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09039_ _05082_ _05084_ _05098_ net593 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[14\]
+ sky130_fd_sc_hd__o32a_4
XFILLER_0_103_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08313__B net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12050_ _07378_ _07468_ _07846_ _07861_ vssd1 vssd1 vccd1 vccd1 _07862_ sky130_fd_sc_hd__o31ai_2
XANTENNA__09357__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold370 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[57\] vssd1 vssd1
+ vccd1 vccd1 net1784 sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[62\] vssd1 vssd1
+ vccd1 vccd1 net1795 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout870_X net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold392 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[33\] vssd1 vssd1
+ vccd1 vccd1 net1806 sky130_fd_sc_hd__dlygate4sd3_1
X_11001_ _06820_ _06821_ vssd1 vssd1 vccd1 vccd1 _06978_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout968_X net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08565__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13646__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12550__S _03678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14331__A team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10372__B1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout850 _04370_ vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__buf_2
Xfanout861 _04296_ vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__buf_2
Xfanout872 net873 vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__buf_2
Xfanout883 net885 vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__clkbuf_2
Xfanout894 _04279_ vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__clkbuf_2
X_15740_ net1307 vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_161_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12952_ net299 net2700 net469 vssd1 vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__mux2_1
Xhold1070 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net2484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net2495 sky130_fd_sc_hd__dlygate4sd3_1
X_11903_ _07597_ _07678_ _07680_ vssd1 vssd1 vccd1 vccd1 _07715_ sky130_fd_sc_hd__and3_1
Xhold1092 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2506 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15671_ net1259 vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_29_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ net287 net2854 net476 vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13381__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17410_ clknet_leaf_65_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[10\]
+ _01106_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15162__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14622_ net1054 vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18390_ net914 vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__clkbuf_1
X_11834_ _07615_ _07617_ _07640_ vssd1 vssd1 vccd1 vccd1 _07646_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09278__D1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09817__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17341_ clknet_leaf_39_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[5\]
+ _01037_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14553_ net1052 vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__inv_2
X_11765_ _07569_ _07571_ _07575_ _07561_ _07547_ vssd1 vssd1 vccd1 vccd1 _07577_ sky130_fd_sc_hd__a311o_1
Xclkbuf_leaf_82_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08096__A2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08047__Y _00040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10978__A2 _06481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10716_ _06709_ _06716_ _04275_ vssd1 vssd1 vccd1 vccd1 _06717_ sky130_fd_sc_hd__o21a_1
X_13504_ net2862 net246 net405 vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__mux2_1
X_17272_ clknet_leaf_30_wb_clk_i _02902_ _00968_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11696_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[16\] team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[17\]
+ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[18\] team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[22\]
+ net994 vssd1 vssd1 vccd1 vccd1 _07508_ sky130_fd_sc_hd__o41a_1
X_14484_ net1068 vssd1 vssd1 vccd1 vccd1 _00114_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_11_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16223_ net1199 vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__inv_2
XANTENNA__08207__C net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13916__A2 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10647_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[6\] team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[5\]
+ _06086_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[7\] vssd1 vssd1
+ vccd1 vccd1 _06652_ sky130_fd_sc_hd__a31o_1
X_13435_ net1995 net234 net414 vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16154_ net1253 vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__inv_2
X_13366_ net2023 net222 net421 vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__mux2_1
X_10578_ net898 _06091_ _06586_ net902 _04175_ vssd1 vssd1 vccd1 vccd1 _06587_ sky130_fd_sc_hd__o32a_1
XFILLER_0_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15105_ net1229 vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__inv_2
X_12317_ _03608_ _03611_ vssd1 vssd1 vccd1 vccd1 _03612_ sky130_fd_sc_hd__or2_2
X_16085_ net1308 vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13297_ net1980 net196 net429 vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__mux2_1
XANTENNA__08223__B net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09348__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12248_ _08010_ _08021_ _03514_ vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__a21oi_1
X_15036_ net1083 vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__inv_2
XANTENNA__12352__A1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[23\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13556__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15337__A net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12460__S net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12179_ _07938_ _07941_ vssd1 vssd1 vccd1 vccd1 _07991_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10363__B1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16987_ clknet_leaf_190_wb_clk_i _02617_ _00683_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15938_ net1289 vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09520__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15869_ net1269 vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__inv_2
XANTENNA__10768__X _06766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13291__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08410_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[29\]
+ net718 _04484_ _04489_ vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__o22a_2
X_17608_ clknet_leaf_81_wb_clk_i _02979_ _01304_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_09390_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[6\]
+ net684 net653 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[6\]
+ _05434_ vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__a221o_1
XANTENNA__08238__X _04321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10487__Y _06500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10418__A1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08341_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[31\]
+ net739 net734 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[31\]
+ _04420_ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__a221o_1
X_17539_ clknet_leaf_81_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[10\]
+ _01235_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11615__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08272_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[14\] _04354_
+ vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08492__C1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_17_Left_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12635__S _03682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09587__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08795__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09339__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08547__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13466__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout496_A net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12370__S net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10354__B1 _06125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11697__A3 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[23\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input1_A ACK_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11494__B net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09726_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[0\]
+ net815 net787 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_87_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09511__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout830_A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout451_X net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09657_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[1\]
+ net756 _05673_ _05677_ _05683_ vssd1 vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout549_X net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout928_A net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08608_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[24\]
+ net709 net657 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__a22o_1
X_09588_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[2\]
+ net774 _05608_ _05614_ _05615_ vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_166_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08539_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[26\]
+ net820 net808 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[26\]
+ _04614_ vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08078__A2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[22\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout716_X net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08308__B net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11550_ _07396_ _07409_ _07412_ _07416_ vssd1 vssd1 vccd1 vccd1 _07461_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_61_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10501_ _06512_ _06513_ net538 vssd1 vssd1 vccd1 vccd1 _06514_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11481_ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[8\] _07391_ net1002
+ vssd1 vssd1 vccd1 vccd1 _07392_ sky130_fd_sc_hd__mux2_1
XANTENNA__12545__S net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13220_ net317 net2506 net350 vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__mux2_1
X_10432_ _06410_ _06447_ net518 vssd1 vssd1 vccd1 vccd1 _06448_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_150_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13151_ net297 net2091 net446 vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__mux2_1
X_10363_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[22\] net904 net536
+ _06380_ vssd1 vssd1 vccd1 vccd1 _06383_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_66_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08250__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10593__B1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12102_ net547 _07600_ vssd1 vssd1 vccd1 vccd1 _07914_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_59_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13082_ net292 net2491 net452 vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__mux2_1
XANTENNA__14323__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input57_A wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10294_ _06312_ _06316_ vssd1 vssd1 vccd1 vccd1 _06317_ sky130_fd_sc_hd__or2_2
XANTENNA__08538__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13376__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12033_ _07365_ net919 _07352_ vssd1 vssd1 vccd1 vccd1 _07845_ sky130_fd_sc_hd__o21ai_1
X_16910_ clknet_leaf_172_wb_clk_i _02540_ _00606_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13229__X _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17890_ clknet_leaf_97_wb_clk_i _03233_ _01586_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16841_ clknet_leaf_25_wb_clk_i _02471_ _00537_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_109_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout680 _04301_ vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__clkbuf_8
Xfanout691 net694 vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__clkbuf_8
X_16772_ clknet_leaf_180_wb_clk_i _02402_ _00468_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13984_ _03834_ _03854_ vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__and2b_1
X_15723_ net1140 vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_126_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09502__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12935_ net243 net2587 net470 vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08710__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15654_ net1249 vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__inv_2
XANTENNA__09602__B net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12866_ net222 net2288 net477 vssd1 vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14605_ net1087 vssd1 vssd1 vccd1 vccd1 _00235_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18373_ net1358 vssd1 vssd1 vccd1 vccd1 la_data_out[21] sky130_fd_sc_hd__buf_2
X_11817_ _07615_ _07617_ vssd1 vssd1 vccd1 vccd1 _07629_ sky130_fd_sc_hd__nand2_1
X_15585_ net1251 vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ net195 net2701 net487 vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_174_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08218__B net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17324_ clknet_leaf_4_wb_clk_i _02954_ _01020_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_174_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14536_ net1223 vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__inv_2
X_11748_ _07531_ _07558_ vssd1 vssd1 vccd1 vccd1 _07560_ sky130_fd_sc_hd__or2_1
XFILLER_0_126_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17255_ clknet_leaf_201_wb_clk_i _02885_ _00951_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12455__S net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14467_ net1203 vssd1 vssd1 vccd1 vccd1 _00097_ sky130_fd_sc_hd__inv_2
X_11679_ _07480_ _07492_ _07493_ net1469 vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__o22a_1
X_16206_ net1281 vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13418_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[8\]
+ net296 net419 vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__mux2_1
X_17186_ clknet_leaf_4_wb_clk_i _02816_ _00882_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_14398_ net1515 vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08777__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16137_ net1274 vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__inv_2
XANTENNA__08241__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13349_ net290 net2939 net424 vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10584__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16068_ net1260 vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__inv_2
XANTENNA__08529__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13286__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15019_ net1070 vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__inv_2
X_08890_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[17\]
+ net836 net751 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10639__A1 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09511_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[4\]
+ net717 _05546_ _05549_ vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_79_748 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11300__A2 _07096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08701__B1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09442_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[17\] net966
+ vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09373_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[7\]
+ net592 _05412_ _05418_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[7\]
+ sky130_fd_sc_hd__o22a_4
XFILLER_0_46_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout244_A net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_25_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08324_ net942 net1014 net925 vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__and3_4
X_08255_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[31\]
+ net677 net626 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[31\]
+ _04326_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__a221o_1
XFILLER_0_89_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_946 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08480__A2 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout411_A _03728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1153_A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08186_ _04267_ _04268_ vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__or2_4
XFILLER_0_132_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10575__B1 _06263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout780_A net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12316__A1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[17\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13196__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout499_X net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09193__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout666_X net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08940__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09703__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09709_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[0\]
+ net951 net937 net926 vssd1 vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__and4_1
X_10981_ _06808_ _06809_ _06864_ net1043 vssd1 vssd1 vccd1 vccd1 _06962_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout833_X net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11444__S net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12720_ net328 net2925 net497 vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12651_ _03686_ _03688_ _07349_ _07351_ vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_100_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11055__A1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11602_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[22\] net993 vssd1
+ vssd1 vccd1 vccd1 _07474_ sky130_fd_sc_hd__and2_2
XFILLER_0_66_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12582_ _03651_ net1802 net204 vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__mux2_1
X_15370_ net1121 vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_152_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14321_ net378 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__nor2_1
X_11533_ net1001 _07443_ _07442_ vssd1 vssd1 vccd1 vccd1 _07444_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08471__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17040_ clknet_leaf_124_wb_clk_i _02670_ _00736_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14252_ team_05_WB.instance_to_wrap.total_design.keypad0.counter\[3\] team_05_WB.instance_to_wrap.total_design.keypad0.counter\[5\]
+ team_05_WB.instance_to_wrap.total_design.keypad0.counter\[6\] team_05_WB.instance_to_wrap.total_design.keypad0.counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__or4b_1
X_11464_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[5\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[5\]
+ net1034 vssd1 vssd1 vccd1 vccd1 _07375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire377 _04858_ vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__buf_4
XANTENNA__08759__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10415_ _06263_ _06431_ net371 vssd1 vssd1 vccd1 vccd1 _06432_ sky130_fd_sc_hd__mux2_1
X_13203_ _06384_ net2812 net351 vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__mux2_1
X_14183_ team_05_WB.EN_VAL_REG net913 vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__or2_1
X_11395_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[9\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[8\]
+ _07324_ vssd1 vssd1 vccd1 vccd1 _07326_ sky130_fd_sc_hd__and3_1
XANTENNA__09420__A1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10346_ _06362_ _06366_ _04264_ vssd1 vssd1 vccd1 vccd1 _06367_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_21_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13134_ net241 net2792 net446 vssd1 vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13065_ net219 net2724 net455 vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__mux2_1
X_17942_ clknet_leaf_33_wb_clk_i _03281_ _01638_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10277_ _06298_ _06299_ net371 vssd1 vssd1 vccd1 vccd1 _06300_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14287__C_N _06918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12016_ _07825_ _07826_ _07827_ vssd1 vssd1 vccd1 vccd1 _07828_ sky130_fd_sc_hd__and3_1
X_17873_ clknet_leaf_99_wb_clk_i _03216_ _01569_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08931__B1 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16824_ clknet_leaf_29_wb_clk_i _02454_ _00520_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_124_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16755_ clknet_leaf_164_wb_clk_i _02385_ _00451_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13967_ team_05_WB.instance_to_wrap.CPU_DAT_O\[4\] net546 _07451_ vssd1 vssd1 vccd1
+ vccd1 _03839_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15706_ net1255 vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__inv_2
X_12918_ net296 net2228 net475 vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16686_ clknet_leaf_173_wb_clk_i _02316_ _00382_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13898_ net1573 net981 _03785_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[20\]
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_17_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15637_ net1282 vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12849_ net290 net2566 net480 vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18356_ net1341 vssd1 vssd1 vccd1 vccd1 la_data_out[4] sky130_fd_sc_hd__buf_2
XFILLER_0_56_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15568_ net1282 vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17307_ clknet_leaf_186_wb_clk_i _02937_ _01003_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_14519_ net1101 vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18287_ net1379 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
X_15499_ net1167 vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08462__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08040_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[4\] vssd1
+ vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17238_ clknet_leaf_141_wb_clk_i _02868_ _00934_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold903 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2317 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold914 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net2328 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12913__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17169_ clknet_leaf_122_wb_clk_i _02799_ _00865_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10557__B1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold925 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2339 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold936 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net2350 sky130_fd_sc_hd__dlygate4sd3_1
Xhold947 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net2361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net2372 sky130_fd_sc_hd__dlygate4sd3_1
Xhold969 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2383 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09991_ _06018_ _06019_ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11529__S net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08942_ _04999_ _05001_ _05003_ _05005_ vssd1 vssd1 vccd1 vccd1 _05006_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12214__A _07476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14132__C net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08873_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[17\]
+ net690 net598 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__a22o_1
XANTENNA__08922__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout194_A _06184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15525__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout459_A _03712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09425_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[5\]
+ net693 net662 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[5\]
+ _05467_ vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__a221o_1
XFILLER_0_137_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout626_A net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09356_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[7\]
+ net838 net779 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05402_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_139_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_139_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_142_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08989__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08307_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[31\]
+ net819 net816 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__a22o_1
X_09287_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[8\]
+ net709 net596 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout414_X net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08238_ net881 _04296_ net859 vssd1 vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout995_A _07470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08305__C net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08169_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[8\] team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[7\]
+ _04249_ vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__and3_2
XANTENNA__12823__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10200_ _06119_ _06131_ net516 vssd1 vssd1 vccd1 vccd1 _06226_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11180_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[39\] _07097_
+ _07111_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[111\] vssd1
+ vssd1 vccd1 vccd1 _07146_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_56_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08602__A _04656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout783_X net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10131_ net514 _06158_ vssd1 vssd1 vccd1 vccd1 _06159_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09166__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08321__B net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10062_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[11\] _06090_ vssd1
+ vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_145_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout950_X net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08913__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13654__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14870_ net1096 vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13821_ team_05_WB.instance_to_wrap.total_design.core.data_mem.state\[0\] team_05_WB.instance_to_wrap.total_design.core.data_mem.state\[2\]
+ _04177_ _03748_ vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__and4_2
XFILLER_0_173_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16540_ clknet_leaf_154_wb_clk_i _02170_ _00236_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13752_ _05212_ _06408_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[20\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_134_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10964_ _06944_ _06948_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[19\]
+ net564 vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_70_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12703_ net248 net2200 net497 vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__mux2_1
X_16471_ clknet_leaf_145_wb_clk_i _02101_ _00167_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13683_ net2233 net302 net385 vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__mux2_1
XANTENNA__12794__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[10\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10895_ net960 _05921_ net565 vssd1 vssd1 vccd1 vccd1 _06892_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08692__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18210_ clknet_leaf_42_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[31\]
+ _01905_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_15422_ net1113 vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__inv_2
X_12634_ net1625 _07798_ _03682_ vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__mux2_1
XANTENNA__08336__X _04418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18254__Q team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18141_ clknet_leaf_163_wb_clk_i _03444_ _01837_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_15353_ net1058 vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__inv_2
X_12565_ _03604_ net1833 net207 vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08444__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08055__Y _04175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14304_ net381 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[31\]
+ net380 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[30\] vssd1
+ vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__a22oi_2
X_18072_ clknet_leaf_85_wb_clk_i _00013_ _01768_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11516_ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[14\] _07426_ net1001
+ vssd1 vssd1 vccd1 vccd1 _07427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15284_ net1076 vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__inv_2
X_12496_ net1645 _03604_ _03674_ vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_670 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17023_ clknet_leaf_155_wb_clk_i _02653_ _00719_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14235_ net1777 _04026_ vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__xor2_1
XFILLER_0_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_117_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11447_ net1050 net1049 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[29\]
+ vssd1 vssd1 vccd1 vccd1 _07358_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12733__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11378_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[2\] _07067_
+ net731 vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__mux2_1
XANTENNA_output88_A net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14166_ net2973 net504 net909 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[15\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10329_ _05929_ _06349_ vssd1 vssd1 vccd1 vccd1 _06350_ sky130_fd_sc_hd__xor2_4
X_13117_ net299 net2718 net450 vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14097_ net910 _03963_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[9\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__08231__B net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17925_ clknet_leaf_42_wb_clk_i _03264_ _01621_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13048_ net280 net2317 net457 vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__mux2_1
Xfanout1250 net1251 vssd1 vssd1 vccd1 vccd1 net1250 sky130_fd_sc_hd__buf_4
XANTENNA__13564__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1261 net1279 vssd1 vssd1 vccd1 vccd1 net1261 sky130_fd_sc_hd__clkbuf_2
X_17856_ clknet_leaf_93_wb_clk_i _03199_ _01552_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[38\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1272 net1278 vssd1 vssd1 vccd1 vccd1 net1272 sky130_fd_sc_hd__buf_4
XANTENNA__13791__C net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1283 net1287 vssd1 vssd1 vccd1 vccd1 net1283 sky130_fd_sc_hd__buf_2
Xfanout1294 net1311 vssd1 vssd1 vccd1 vccd1 net1294 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_1_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12688__B net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11592__B _07472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16807_ clknet_leaf_199_wb_clk_i _02437_ _00503_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17787_ clknet_leaf_78_wb_clk_i _03130_ _01483_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[97\]
+ sky130_fd_sc_hd__dfrtp_1
X_14999_ net1096 vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__inv_2
XFILLER_0_163_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16738_ clknet_leaf_7_wb_clk_i _02368_ _00434_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16669_ clknet_leaf_131_wb_clk_i _02299_ _00365_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16176__A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12908__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11019__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15080__A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09210_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[10\]
+ net841 net786 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[10\]
+ _05261_ vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__a221o_1
X_18408_ net914 vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09141_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[11\]
+ net695 net610 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__a22o_1
X_18339_ net1328 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
XFILLER_0_115_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09072_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[13\]
+ net790 net756 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05130_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12519__A1 _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14341__A1_N _05596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12643__S net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold700 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2114 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold711 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold722 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2136 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold733 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 net2147 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09518__A _05556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold744 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 net2158 sky130_fd_sc_hd__dlygate4sd3_1
Xhold755 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2169 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_39_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__17508__Q team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[11\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold766 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2180 sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 net2191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2202 sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ _06002_ _05531_ vssd1 vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__nand2b_4
Xhold799 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2213 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08925_ _04989_ vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_51_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout576_A net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1400 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2814 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13474__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1411 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2825 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1422 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net2836 sky130_fd_sc_hd__dlygate4sd3_1
X_08856_ _04922_ vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__inv_2
Xhold1433 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net2847 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10702__B1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1444 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1455 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1466 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net2880 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1477 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net2891 sky130_fd_sc_hd__dlygate4sd3_1
X_08787_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[19\]
+ net715 _04854_ _04857_ vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_19_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1488 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2902 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout743_A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1499 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 net2913 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09320__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12818__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08674__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout629_X net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Left_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09408_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[6\]
+ net802 net737 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05452_ sky130_fd_sc_hd__a22o_1
X_10680_ _06398_ _06508_ _06545_ net332 _06681_ vssd1 vssd1 vccd1 vccd1 _06683_ sky130_fd_sc_hd__o221a_1
XANTENNA__09700__B _05731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09339_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[7\]
+ net708 net622 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05386_ sky130_fd_sc_hd__a22o_1
XANTENNA__08426__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11023__A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_78_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_63_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12350_ net545 _07476_ net354 vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__o21a_2
XFILLER_0_50_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11301_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[9\] _07101_ _07108_
+ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[89\] vssd1 vssd1 vccd1
+ vccd1 _07261_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13649__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12281_ _03575_ _07986_ vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__and2b_1
XANTENNA__12553__S net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14020_ _03887_ _03889_ vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__nor2_1
X_11232_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[44\] _07091_
+ _07097_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[36\] vssd1 vssd1
+ vccd1 vccd1 _07195_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09387__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11194__B1 _07110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11163_ _07087_ _07078_ _07059_ vssd1 vssd1 vccd1 vccd1 _07129_ sky130_fd_sc_hd__and3b_4
XTAP_TAPCELL_ROW_112_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_36_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_8_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10941__B1 _06898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09139__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10114_ net376 net367 vssd1 vssd1 vccd1 vccd1 _06142_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_164_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11094_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[2\] _07033_
+ vssd1 vssd1 vccd1 vccd1 _07061_ sky130_fd_sc_hd__nand2_1
X_15971_ net1304 vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_164_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17710_ clknet_leaf_87_wb_clk_i _03053_ _01406_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[84\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13384__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14922_ net1109 vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__inv_2
X_10045_ _04573_ net363 vssd1 vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold60 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[0\]
+ vssd1 vssd1 vccd1 vccd1 net1474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[21\]
+ vssd1 vssd1 vccd1 vccd1 net1485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[18\] vssd1 vssd1
+ vccd1 vccd1 net1496 sky130_fd_sc_hd__dlygate4sd3_1
X_17641_ clknet_leaf_68_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[8\]
+ _01337_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_14853_ net1203 vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__inv_2
Xhold93 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[8\]
+ vssd1 vssd1 vccd1 vccd1 net1507 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_output126_A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13804_ net1600 net971 net724 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[15\]
+ sky130_fd_sc_hd__and3_1
X_17572_ clknet_leaf_110_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[9\]
+ _01268_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_14784_ net1199 vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__inv_2
XANTENNA__10102__A net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08114__A1 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11996_ _07803_ _07805_ _07806_ _07807_ vssd1 vssd1 vccd1 vccd1 _07808_ sky130_fd_sc_hd__or4_1
XANTENNA__12020__C _07821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09311__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16523_ clknet_leaf_188_wb_clk_i _02153_ _00219_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13735_ net922 _06706_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[3\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_133_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10947_ _06934_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[22\] net564
+ vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__mux2_1
XANTENNA__12728__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08665__A2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16454_ clknet_leaf_116_wb_clk_i _02084_ _00150_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13666_ net2217 net234 net385 vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__mux2_1
X_10878_ _06796_ _06874_ _06793_ _06794_ vssd1 vssd1 vccd1 vccd1 _06875_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_119_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10756__B _05801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15405_ net1131 vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12617_ net1620 _07789_ _03682_ vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_119_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16385_ clknet_leaf_148_wb_clk_i _02015_ _00081_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08417__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13597_ net2775 net222 net394 vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08226__B net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18124_ clknet_leaf_48_wb_clk_i _00038_ _01820_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15336_ net1219 vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__inv_2
X_12548_ _03651_ net1872 net205 vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09090__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18055_ net1037 _03393_ _01751_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_41_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12463__S _03670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15267_ net1206 vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__inv_2
X_12479_ net1749 _03651_ net211 vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__mux2_1
XANTENNA_2 _06518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17006_ clknet_leaf_170_wb_clk_i _02636_ _00702_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_14218_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[13\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[12\]
+ _04011_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[14\] vssd1
+ vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__a31o_1
XANTENNA_wire377_A _04858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15198_ net1056 vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__inv_2
XANTENNA__11185__B1 _07118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14149_ team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.next_next_data_read
+ team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.next_next_fetch _03684_ vssd1
+ vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__and3b_1
Xfanout509 _07295_ vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__buf_2
XFILLER_0_120_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13294__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08710_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[22\]
+ net848 net750 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__a22o_1
X_17908_ clknet_leaf_77_wb_clk_i _03251_ _01604_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_09690_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[1\]
+ net665 _05707_ _05708_ _05710_ vssd1 vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__a2111o_1
Xfanout1080 net1086 vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__buf_2
XANTENNA__09550__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1091 net1094 vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__buf_4
X_08641_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[24\]
+ net592 _04709_ _04715_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[24\]
+ sky130_fd_sc_hd__o22a_4
XFILLER_0_174_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17839_ clknet_leaf_87_wb_clk_i _03182_ _01535_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[85\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12211__B net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12437__A0 _03623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08572_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[25\]
+ net650 net627 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[25\]
+ _04647_ vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__a221o_1
XANTENNA__10012__A net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09801__A _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12638__S net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08656__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_112_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14419__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08408__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09124_ _05173_ _05175_ _05177_ _05179_ vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__or4_1
XFILLER_0_44_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09081__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13469__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09055_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[13\]
+ net690 net644 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__a22o_1
XANTENNA__12373__S _07852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1233_A net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09369__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold530 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net1944 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08152__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11176__B1 _07123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout693_A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold541 net118 vssd1 vssd1 vccd1 vccd1 net1955 sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 _07334_ vssd1 vssd1 vccd1 vccd1 net1966 sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 net97 vssd1 vssd1 vccd1 vccd1 net1977 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold574 net102 vssd1 vssd1 vccd1 vccd1 net1988 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1021_X net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold585 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net1999 sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net2010 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09957_ _04778_ _04797_ vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout481_X net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout860_A net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout958_A net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08908_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[16\]
+ net699 net632 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[16\]
+ _04971_ vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__a221o_1
XANTENNA__09254__Y _05305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09888_ _04594_ _05912_ _05916_ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_151_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold1230 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 net2644 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09541__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1241 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2655 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1252 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2666 sky130_fd_sc_hd__dlygate4sd3_1
X_08839_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[18\]
+ net822 net737 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__a22o_1
XANTENNA__13217__B net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1263 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2677 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1274 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net2688 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout746_X net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08895__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1285 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2699 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15713__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1296 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2710 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11850_ _07656_ _07659_ _07653_ _07654_ vssd1 vssd1 vccd1 vccd1 _07662_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_68_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_154_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_154_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10801_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[20\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[20\]
+ vssd1 vssd1 vccd1 vccd1 _06798_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_68_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12548__S net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08647__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11781_ _07591_ _07592_ vssd1 vssd1 vccd1 vccd1 _07593_ sky130_fd_sc_hd__nor2_1
XANTENNA__11452__S net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11305__X _07265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13520_ net2015 net313 net406 vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__mux2_1
X_10732_ net334 _06277_ _06730_ net554 _06722_ vssd1 vssd1 vccd1 vccd1 _06732_ sky130_fd_sc_hd__o221a_1
XFILLER_0_83_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13451_ net2900 net296 net415 vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__mux2_1
X_10663_ net333 _06125_ _06503_ _06526_ _06666_ vssd1 vssd1 vccd1 vccd1 _06667_ sky130_fd_sc_hd__o221a_1
XFILLER_0_137_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12402_ net1900 _03641_ net216 vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__mux2_1
X_16170_ net1143 vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10594_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[9\] _06089_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06602_ sky130_fd_sc_hd__a21oi_1
X_13382_ net2316 net292 net420 vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__mux2_1
XANTENNA__09072__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15121_ net1188 vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__inv_2
XANTENNA__13379__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12333_ net354 _03599_ _03626_ _03616_ _07506_ vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_114_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09158__A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15052_ net1109 vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__inv_2
X_12264_ _07968_ _07977_ _03558_ vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__and3_1
XANTENNA__11167__B1 _07110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_190_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14003_ _03872_ _03873_ vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__and2b_1
X_11215_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[125\] _07099_
+ _07126_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[85\] _07178_
+ vssd1 vssd1 vccd1 vccd1 _07179_ sky130_fd_sc_hd__a221o_1
X_12195_ _08006_ vssd1 vssd1 vccd1 vccd1 _08007_ sky130_fd_sc_hd__inv_2
XANTENNA__08997__A _05034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__clkbuf_4
X_11146_ _07039_ _07088_ vssd1 vssd1 vccd1 vccd1 _07112_ sky130_fd_sc_hd__or2_4
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 ADR_O[27] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11077_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[2\] team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[1\]
+ vssd1 vssd1 vccd1 vccd1 _07044_ sky130_fd_sc_hd__nand2_1
X_15954_ net1289 vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__inv_2
XANTENNA__12312__A _03604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10028_ _04157_ _06054_ vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__nand2_1
XANTENNA__09532__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14905_ net1051 vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__inv_2
X_15885_ net1269 vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__inv_2
XANTENNA__12419__A0 _03614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17624_ clknet_leaf_66_wb_clk_i _02995_ _01320_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_14836_ net1068 vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17555_ clknet_leaf_62_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[26\]
+ _01251_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12458__S _03670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14767_ net1280 vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__inv_2
XANTENNA__10767__A net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11979_ _07790_ _07787_ _07518_ _07512_ vssd1 vssd1 vccd1 vccd1 _07791_ sky130_fd_sc_hd__o2bb2a_4
XANTENNA__08638__A2 _04366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16506_ clknet_leaf_10_wb_clk_i _02136_ _00202_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13718_ net905 _06445_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[18\]
+ sky130_fd_sc_hd__and2_1
X_17486_ clknet_leaf_36_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[21\]
+ _01182_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14698_ net1110 vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13919__B1 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16437_ clknet_leaf_22_wb_clk_i _02067_ _00133_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13649_ net2845 net295 net391 vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__mux2_1
XANTENNA__09599__B1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16368_ clknet_leaf_152_wb_clk_i _01998_ _00064_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18107_ clknet_leaf_54_wb_clk_i _03430_ _01803_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[24\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_42_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13289__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15319_ net1096 vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16299_ net1154 vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18038_ clknet_leaf_94_wb_clk_i _03376_ _01734_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12921__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout306 net308 vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__buf_1
X_09811_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[20\]
+ net682 net629 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__a22o_1
Xfanout317 _06671_ vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__clkbuf_2
Xfanout328 _06705_ vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__clkbuf_2
Xfanout339 _03693_ vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__buf_4
XFILLER_0_158_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09742_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[0\]
+ net887 _04287_ net866 vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__and4_1
XANTENNA__12222__A _07774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14140__C net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09523__B1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09673_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[1\]
+ net883 net871 net857 vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__and4_1
XANTENNA__08877__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08624_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[24\]
+ net788 net776 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__a22o_1
XANTENNA__10684__A2 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08555_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[26\]
+ net593 _04627_ _04631_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[26\]
+ sky130_fd_sc_hd__o22a_2
XANTENNA__12368__S net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17521__Q team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[24\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08629__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout441_A _03716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1183_A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout539_A net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08486_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[27\]
+ net688 net657 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout706_A _04292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout327_X net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_99_Left_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09054__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09107_ _05150_ _05151_ _05162_ _05163_ vssd1 vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__or4_1
XANTENNA__13199__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08801__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14335__B1 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09038_ _05086_ _05091_ _05093_ _05097_ vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout696_X net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08313__C net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold360 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[85\] vssd1 vssd1
+ vccd1 vccd1 net1774 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12831__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold371 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[76\] vssd1 vssd1
+ vccd1 vccd1 net1785 sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[54\] vssd1 vssd1
+ vccd1 vccd1 net1796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[88\] vssd1 vssd1
+ vccd1 vccd1 net1807 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ _06977_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[12\] net568
+ vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__mux2_1
XANTENNA__10372__A1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout863_X net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout840 _04377_ vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__buf_4
Xfanout851 _04370_ vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__clkbuf_8
Xfanout862 net863 vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__buf_2
XANTENNA__11674__C net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout873 _04284_ vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__clkbuf_2
Xfanout884 net885 vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__clkbuf_2
Xfanout895 net898 vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12951_ net286 net2859 net468 vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__mux2_1
Xhold1060 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[11\] vssd1 vssd1
+ vccd1 vccd1 net2474 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11321__B1 _07102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08868__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1071 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2485 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13662__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11902_ _07529_ _07713_ vssd1 vssd1 vccd1 vccd1 _07714_ sky130_fd_sc_hd__nor2_1
X_15670_ net1256 vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__inv_2
Xhold1082 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2496 sky130_fd_sc_hd__dlygate4sd3_1
X_12882_ net290 net2833 net476 vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__mux2_1
Xhold1093 net134 vssd1 vssd1 vccd1 vccd1 net2507 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09441__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[25\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14621_ net1090 vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__inv_2
X_11833_ _07629_ _07640_ _07642_ _07638_ vssd1 vssd1 vccd1 vccd1 _07645_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_159_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17340_ clknet_leaf_41_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[4\]
+ _01036_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14552_ net1242 vssd1 vssd1 vccd1 vccd1 _00182_ sky130_fd_sc_hd__inv_2
XANTENNA__11624__B2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11764_ _07572_ _07575_ _07562_ vssd1 vssd1 vccd1 vccd1 _07576_ sky130_fd_sc_hd__a21boi_1
XPHY_EDGE_ROW_161_Right_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09293__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13503_ net2523 net226 net406 vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_155_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10715_ _06432_ net347 _06715_ vssd1 vssd1 vccd1 vccd1 _06716_ sky130_fd_sc_hd__o21ai_1
X_17271_ clknet_leaf_144_wb_clk_i _02901_ _00967_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_155_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14483_ net1213 vssd1 vssd1 vccd1 vccd1 _00113_ sky130_fd_sc_hd__inv_2
X_11695_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[29\] net995 vssd1
+ vssd1 vccd1 vccd1 _07507_ sky130_fd_sc_hd__and2_1
X_16222_ net1181 vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__inv_2
X_13434_ net2132 net241 net414 vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__mux2_1
X_10646_ _06642_ _06649_ _06650_ net538 vssd1 vssd1 vccd1 vccd1 _06651_ sky130_fd_sc_hd__a31o_1
XFILLER_0_64_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16153_ net1255 vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__inv_2
XANTENNA__08253__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10526__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13365_ net1964 net220 net422 vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_51_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10577_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[11\] _06090_ vssd1
+ vssd1 vccd1 vccd1 _06586_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15104_ net1199 vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__inv_2
X_12316_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[17\] net1000 _03511_
+ _03589_ net544 vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__a221o_1
XANTENNA__14326__B1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[12\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16084_ net1308 vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__inv_2
X_13296_ net2112 net198 net429 vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08223__C net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15035_ net1098 vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__inv_2
X_12247_ _03517_ _03531_ _03536_ _03540_ vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__nor4_1
XANTENNA__12741__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08556__A1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12352__A2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[30\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12178_ _07988_ _07989_ vssd1 vssd1 vccd1 vccd1 _07990_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10363__B2 _06380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11129_ _07078_ _07093_ vssd1 vssd1 vccd1 vccd1 _07095_ sky130_fd_sc_hd__nand2_2
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16986_ clknet_leaf_31_wb_clk_i _02616_ _00682_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09505__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15937_ net1271 vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__inv_2
XANTENNA__11312__B1 _07121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08859__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13572__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15868_ net1310 vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__inv_2
X_17607_ clknet_leaf_81_wb_clk_i _02978_ _01303_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_14819_ net1207 vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__inv_2
X_15799_ net1302 vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11615__A1 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08340_ net942 net938 _04418_ vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__and3_1
XFILLER_0_171_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17538_ clknet_leaf_81_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[9\]
+ _01234_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11615__B2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09284__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08271_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[13\] net1019
+ _04353_ vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__or3b_1
XFILLER_0_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17469_ clknet_leaf_40_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[4\]
+ _01165_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__12916__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13160__X _03716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09036__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08244__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14135__C net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14317__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17516__Q team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[19\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout391_A _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10354__B2 _06355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11697__A4 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[30\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout489_A _03700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14096__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09725_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[0\]
+ net837 net781 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_87_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout656_A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13482__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09656_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[1\]
+ net821 _05679_ _05682_ _05684_ vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_59_1092 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08607_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[24\]
+ net714 net600 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[24\]
+ _04681_ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout823_A net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09587_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[2\]
+ net770 _05603_ _05607_ _05620_ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout444_X net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1186_X net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08538_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[26\]
+ net839 net766 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11606__B2 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[19\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09275__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_102_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08308__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08483__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12826__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout611_X net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08469_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[28\]
+ net852 net848 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[28\]
+ _04547_ vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__a221o_1
XFILLER_0_108_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout709_X net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10500_ _06033_ _06049_ _06502_ net554 vssd1 vssd1 vccd1 vccd1 _06513_ sky130_fd_sc_hd__o22a_1
XFILLER_0_80_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11480_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[8\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[8\]
+ net1034 vssd1 vssd1 vccd1 vccd1 _07391_ sky130_fd_sc_hd__mux2_1
XANTENNA__09027__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10431_ _06142_ _06153_ vssd1 vssd1 vccd1 vccd1 _06447_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_150_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08324__B net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13150_ net298 net2226 net445 vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__mux2_1
X_10362_ _06098_ _06381_ vssd1 vssd1 vccd1 vccd1 _06382_ sky130_fd_sc_hd__or2_2
XFILLER_0_104_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13657__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12101_ _07864_ _07902_ _07910_ vssd1 vssd1 vccd1 vccd1 _07913_ sky130_fd_sc_hd__nand3_1
XFILLER_0_130_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12561__S net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10293_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[25\] net904 net968
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[25\] _06315_ vssd1
+ vssd1 vccd1 vccd1 _06316_ sky130_fd_sc_hd__a221o_1
X_13081_ net280 net2290 net453 vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__mux2_1
XANTENNA__14342__A _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12032_ _07363_ _07843_ vssd1 vssd1 vccd1 vccd1 _07844_ sky130_fd_sc_hd__nor2_1
Xhold190 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[75\] vssd1 vssd1
+ vccd1 vccd1 net1604 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10345__A1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16840_ clknet_leaf_197_wb_clk_i _02470_ _00536_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_109_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout670 net671 vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__buf_4
Xfanout681 _04301_ vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__buf_4
X_16771_ clknet_leaf_192_wb_clk_i _02401_ _00467_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout692 net694 vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__clkbuf_8
X_13983_ _03852_ _03853_ _03834_ vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__and3b_1
XANTENNA__12098__B2 _07864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13392__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15722_ net1142 vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_126_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12934_ net223 net2208 net469 vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08339__X _04421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18257__Q team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[11\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15653_ net1249 vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__inv_2
X_12865_ net218 net2151 net478 vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__mux2_1
XANTENNA__09602__C net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ net1109 vssd1 vssd1 vccd1 vccd1 _00234_ sky130_fd_sc_hd__inv_2
X_18372_ net1357 vssd1 vssd1 vccd1 vccd1 la_data_out[20] sky130_fd_sc_hd__buf_2
X_11816_ _07621_ _07625_ _07627_ vssd1 vssd1 vccd1 vccd1 _07628_ sky130_fd_sc_hd__a21oi_4
X_15584_ net1251 vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__inv_2
XANTENNA__09266__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12796_ net197 net2231 net487 vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_174_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ clknet_leaf_162_wb_clk_i _02953_ _01019_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[19\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_174_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ net1199 vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_174_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11747_ _07548_ _07558_ _07531_ vssd1 vssd1 vccd1 vccd1 _07559_ sky130_fd_sc_hd__o21ba_1
XANTENNA__12736__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17254_ clknet_leaf_115_wb_clk_i _02884_ _00950_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10281__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14466_ net1217 vssd1 vssd1 vccd1 vccd1 _00096_ sky130_fd_sc_hd__inv_2
X_11678_ team_05_WB.instance_to_wrap.wishbone.curr_state\[0\] _07344_ _07491_ vssd1
+ vssd1 vccd1 vccd1 _07493_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16205_ net1184 vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13417_ net2636 net301 net418 vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10629_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[8\] _06088_ vssd1
+ vssd1 vccd1 vccd1 _06635_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17185_ clknet_leaf_147_wb_clk_i _02815_ _00881_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_14397_ net1511 vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08234__B net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16136_ net1273 vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13348_ net278 net2918 net424 vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13567__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16067_ net1260 vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__inv_2
XANTENNA__12471__S net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13794__C net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13279_ net270 net2618 net432 vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15018_ net1109 vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__inv_2
XANTENNA__09726__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16969_ clknet_leaf_20_wb_clk_i _02599_ _00665_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16179__A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09510_ _05533_ _05536_ _05538_ _05548_ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__or4_1
XFILLER_0_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09441_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[25\] _05306_
+ vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18394__A net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09372_ _05414_ _05415_ _05416_ _05417_ vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08323_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[31\]
+ net779 net775 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[31\]
+ _04402_ vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__a221o_1
XANTENNA__08465__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09662__C1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout237_A _06346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08254_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[31\]
+ net608 _04336_ net721 vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__a211o_1
XANTENNA__09009__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10674__B net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12013__A1 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[30\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08185_ _04231_ _04241_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__nor2_4
XFILLER_0_104_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout404_A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1146_A net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_502 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10024__B1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11221__C1 _07031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13477__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12381__S net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout394_X net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout773_A _04406_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13277__A0 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout561_X net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout659_X net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09708_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[0\]
+ net944 net936 net929 vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__and4_1
X_10980_ _06808_ _06809_ _06864_ vssd1 vssd1 vccd1 vccd1 _06961_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09496__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09639_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[1\]
+ net948 net935 net925 vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__and4_1
XANTENNA__13225__B net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout826_X net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08319__B net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12650_ team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.state\[0\] team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.state\[2\]
+ team_05_WB.instance_to_wrap.total_design.core.mem_ctrl.state\[1\] vssd1 vssd1 vccd1
+ vccd1 _03688_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_168_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09248__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11601_ net123 net1011 net346 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__a22o_1
XANTENNA__12556__S net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12581_ _03662_ net1852 net204 vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__mux2_1
XANTENNA__08456__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11460__S net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14320_ _05035_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__nor2_1
X_11532_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[13\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[13\]
+ net1033 vssd1 vssd1 vccd1 vccd1 _07443_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08335__A net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14251_ team_05_WB.instance_to_wrap.total_design.keypad0.counter\[4\] _04018_ vssd1
+ vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__xor2_1
XFILLER_0_151_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11463_ net920 _07371_ _07373_ vssd1 vssd1 vccd1 vccd1 _07374_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13202_ net230 net2682 net352 vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__mux2_1
Xwire378 _04736_ vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__buf_4
XFILLER_0_21_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10414_ _06358_ _06430_ net528 vssd1 vssd1 vccd1 vccd1 _06431_ sky130_fd_sc_hd__mux2_1
X_14182_ net1609 net506 net909 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[31\]
+ sky130_fd_sc_hd__and3_1
X_11394_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[8\] _07324_
+ vssd1 vssd1 vccd1 vccd1 _07325_ sky130_fd_sc_hd__and2_1
XANTENNA__09420__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13387__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13133_ net243 net2205 net446 vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__mux2_1
X_10345_ net895 _06364_ _06365_ vssd1 vssd1 vccd1 vccd1 _06366_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_104_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17941_ clknet_leaf_35_wb_clk_i _03280_ _01637_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13064_ net191 net2891 net455 vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10276_ _06206_ _06208_ net526 vssd1 vssd1 vccd1 vccd1 _06299_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_167_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12015_ _07478_ _07507_ _07523_ _07601_ _07449_ vssd1 vssd1 vccd1 vccd1 _07827_ sky130_fd_sc_hd__a41o_1
X_17872_ clknet_leaf_104_wb_clk_i _03215_ _01568_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10105__A _05078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16823_ clknet_leaf_146_wb_clk_i _02453_ _00519_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13966_ net910 _03838_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[3\]
+ sky130_fd_sc_hd__nor2_1
X_16754_ clknet_leaf_123_wb_clk_i _02384_ _00450_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09487__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15705_ net1255 vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__inv_2
X_12917_ net299 net2485 net474 vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__mux2_1
XANTENNA__12491__A1 _03632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11294__A2 _07097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16685_ clknet_leaf_161_wb_clk_i _02315_ _00381_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08695__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13897_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[20\]
+ net558 net574 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[20\]
+ net985 vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_17_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08229__B net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12848_ net280 net2790 net480 vssd1 vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__mux2_1
X_15636_ net1280 vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09239__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_730 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12466__S net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18355_ net1340 vssd1 vssd1 vccd1 vccd1 la_data_out[3] sky130_fd_sc_hd__buf_2
XANTENNA__08447__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15567_ net1246 vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__inv_2
XANTENNA__12319__X _03614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12779_ net282 net2894 net489 vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__mux2_1
XANTENNA__11370__S _06769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14518_ net1084 vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__inv_2
X_17306_ clknet_leaf_13_wb_clk_i _02936_ _01002_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_15498_ net1161 vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18286_ net1378 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
XFILLER_0_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14449_ net1188 vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17237_ clknet_leaf_21_wb_clk_i _02867_ _00933_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17168_ clknet_leaf_152_wb_clk_i _02798_ _00864_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold904 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net2318 sky130_fd_sc_hd__dlygate4sd3_1
Xhold915 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2329 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09411__A2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold926 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2340 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13297__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16119_ net1134 vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__inv_2
Xhold937 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2351 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_29_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold948 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2362 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold959 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2373 sky130_fd_sc_hd__dlygate4sd3_1
X_17099_ clknet_leaf_189_wb_clk_i _02729_ _00795_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_09990_ _05256_ net366 vssd1 vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__or2_1
X_08941_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[16\]
+ net818 net790 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[16\]
+ _05004_ vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_0_wb_clk_i_A wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08872_ _04933_ _04934_ _04936_ _04938_ vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_32_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08383__C1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09478__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12482__A1 _03657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08686__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09424_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[5\]
+ net696 net600 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05467_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09355_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[7\]
+ net827 net747 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__a22o_1
XANTENNA__08438__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12376__S net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10685__A _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout521_A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout619_A net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10245__B1 _06267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08306_ net1016 net942 net928 vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__and3_4
XANTENNA__11588__A3 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_68_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09286_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[8\]
+ net619 net616 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08237_ net879 net874 net860 vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__and3_4
XFILLER_0_132_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout407_X net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_179_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_179_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08168_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[7\] _04249_
+ vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout890_A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09402__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_108_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_108_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_127_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08610__B1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08099_ net1029 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_56_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13000__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10130_ net381 net363 _06157_ vssd1 vssd1 vccd1 vccd1 _06158_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_101_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_128_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout776_X net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10061_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[10\] team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[9\]
+ _06089_ vssd1 vssd1 vccd1 vccd1 _06090_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_73_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11963__B _07774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11455__S net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13820_ net1586 net974 net725 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[31\]
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_162_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09469__A2 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13751_ _05212_ _06424_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[19\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_134_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11276__A2 _07117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10963_ _06898_ _06945_ _06946_ _06947_ vssd1 vssd1 vccd1 vccd1 _06948_ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08677__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13670__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12702_ net226 net2732 net498 vssd1 vssd1 vccd1 vccd1 _02924_ sky130_fd_sc_hd__mux2_1
X_16470_ clknet_leaf_141_wb_clk_i _02100_ _00166_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13682_ net2105 net295 net386 vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__mux2_1
X_10894_ _06888_ _06889_ _06890_ vssd1 vssd1 vccd1 vccd1 _06891_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15421_ net1117 vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__inv_2
X_12633_ _03604_ net1810 net201 vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15352_ net1201 vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__inv_2
X_18140_ clknet_leaf_110_wb_clk_i _03443_ _01836_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_12564_ _03664_ net1800 net205 vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14303_ _04533_ _04552_ vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__nor2_1
X_18071_ clknet_leaf_85_wb_clk_i _00012_ _01767_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11515_ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_i\[14\]
+ team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[14\]
+ net1033 vssd1 vssd1 vccd1 vccd1 _07426_ sky130_fd_sc_hd__mux2_1
X_15283_ net1214 vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12495_ net1726 _03664_ net211 vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17022_ clknet_leaf_163_wb_clk_i _02652_ _00718_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_14234_ _04027_ _04028_ vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_117_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_44_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11446_ net1632 net1007 net727 _07357_ vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18270__Q team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[24\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11200__A2 _07113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14165_ net1906 net502 net908 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[14\]
+ sky130_fd_sc_hd__and3_1
X_11377_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[3\] _07063_
+ net731 vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13116_ net288 net2576 net448 vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__mux2_1
X_10328_ _04798_ _05891_ vssd1 vssd1 vccd1 vccd1 _06349_ sky130_fd_sc_hd__or2_2
X_14096_ net2975 net507 _03962_ vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_147_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08231__C net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17924_ clknet_leaf_43_wb_clk_i _03263_ _01620_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13047_ net285 net2487 net457 vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10259_ _06234_ _06282_ net520 vssd1 vssd1 vccd1 vccd1 _06283_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1240 net1241 vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__clkbuf_4
Xfanout1251 net1252 vssd1 vssd1 vccd1 vccd1 net1251 sky130_fd_sc_hd__buf_4
Xfanout1262 net1264 vssd1 vssd1 vccd1 vccd1 net1262 sky130_fd_sc_hd__buf_4
X_17855_ clknet_leaf_85_wb_clk_i _03198_ _01551_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[37\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1273 net1278 vssd1 vssd1 vccd1 vccd1 net1273 sky130_fd_sc_hd__buf_4
XANTENNA__08380__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_53_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1284 net1285 vssd1 vssd1 vccd1 vccd1 net1284 sky130_fd_sc_hd__buf_4
Xfanout1295 net1298 vssd1 vssd1 vccd1 vccd1 net1295 sky130_fd_sc_hd__buf_4
X_16806_ clknet_leaf_116_wb_clk_i _02436_ _00502_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_17786_ clknet_leaf_91_wb_clk_i _03129_ _01482_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[96\]
+ sky130_fd_sc_hd__dfrtp_1
X_14998_ net1091 vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__inv_2
XANTENNA__12464__A1 _03605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11267__A2 _07091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16737_ clknet_leaf_151_wb_clk_i _02367_ _00433_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08668__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13949_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[6\] team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__or2_1
XFILLER_0_163_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_102_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13580__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16668_ clknet_leaf_157_wb_clk_i _02298_ _00364_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18407_ net1375 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__buf_2
X_15619_ net1173 vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16599_ clknet_leaf_143_wb_clk_i _02229_ _00295_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_09140_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[11\]
+ net711 net598 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[11\]
+ _05194_ vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__a221o_1
X_18338_ net1327 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
XFILLER_0_8_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09093__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_6_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_115_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09071_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[13\]
+ net805 net771 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18269_ clknet_leaf_26_wb_clk_i _03498_ _01964_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08840__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12924__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold701 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net2115 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_201_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_201_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_40_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold712 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net2126 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08199__A2 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold723 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 net2137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold734 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net2148 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold745 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 net2159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold756 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net2170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net2192 sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ _04157_ _04274_ vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__nand2_2
Xhold789 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2203 sky130_fd_sc_hd__dlygate4sd3_1
X_08924_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[16\]
+ net715 _04984_ _04988_ vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__o22a_4
XANTENNA_fanout1011_A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1401 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 net2815 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_141_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1109_A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Left_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1412 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[12\] vssd1 vssd1
+ vccd1 vccd1 net2826 sky130_fd_sc_hd__dlygate4sd3_1
X_08855_ net376 _04921_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__or2_1
Xhold1423 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 net2837 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17524__Q team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[27\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1434 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 net2848 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout569_A _06774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1445 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 net2859 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1456 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2870 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08371__A2 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08786_ _04841_ _04844_ _04846_ _04856_ vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__or4_2
Xhold1467 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 net2881 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1478 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 net2892 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_140_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1489 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2903 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_140_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11258__A2 _07101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12455__A1 _03612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08659__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13490__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09540__Y _05577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09407_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[6\]
+ net827 net742 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[6\]
+ _05450_ vssd1 vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__a221o_1
XFILLER_0_82_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout903_A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09338_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[7\]
+ net653 net603 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[7\]
+ _05383_ vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_80_Left_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09084__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09623__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09269_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[9\]
+ net843 net749 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[9\]
+ _05318_ vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__a221o_1
XANTENNA__12834__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11300_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[89\] _07096_
+ _07129_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[57\] _07247_
+ vssd1 vssd1 vccd1 vccd1 _07260_ sky130_fd_sc_hd__a221o_1
X_12280_ _03573_ _03574_ _03568_ vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__a21boi_2
XTAP_TAPCELL_ROW_75_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11231_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[116\] _07104_
+ _07128_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[68\] _07193_
+ vssd1 vssd1 vccd1 vccd1 _07194_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_180_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08332__B net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08595__C1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11162_ _07038_ _07059_ _07078_ vssd1 vssd1 vccd1 vccd1 _07128_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_112_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13665__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10113_ _06125_ _06140_ net372 vssd1 vssd1 vccd1 vccd1 _06141_ sky130_fd_sc_hd__mux2_1
X_11093_ _07059_ vssd1 vssd1 vccd1 vccd1 _07060_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_164_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15970_ net1288 vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__inv_2
XANTENNA__14350__A _04082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input32_A DAT_I[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ net371 _06048_ vssd1 vssd1 vccd1 vccd1 _06073_ sky130_fd_sc_hd__nand2_1
X_14921_ net1225 vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__inv_2
Xhold50 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[23\] vssd1 vssd1
+ vccd1 vccd1 net1464 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_76_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08362__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold61 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[29\]
+ vssd1 vssd1 vccd1 vccd1 net1475 sky130_fd_sc_hd__dlygate4sd3_1
X_17640_ clknet_leaf_79_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[7\]
+ _01336_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold72 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[14\]
+ vssd1 vssd1 vccd1 vccd1 net1486 sky130_fd_sc_hd__dlygate4sd3_1
X_14852_ net1230 vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__inv_2
Xhold83 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[4\]
+ vssd1 vssd1 vccd1 vccd1 net1497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[14\]
+ vssd1 vssd1 vccd1 vccd1 net1508 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09157__A_N net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13803_ net1575 net970 net723 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[14\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__12446__A1 _07791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11249__A2 _07100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14783_ net1179 vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__inv_2
X_17571_ clknet_leaf_109_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[8\]
+ _01267_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11995_ _07474_ _07518_ _07800_ _07516_ vssd1 vssd1 vccd1 vccd1 _07807_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08114__A2 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13734_ net922 _06729_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[2\]
+ sky130_fd_sc_hd__nor2_1
X_16522_ clknet_leaf_195_wb_clk_i _02152_ _00218_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10946_ net956 _06369_ _06932_ _06933_ vssd1 vssd1 vccd1 vccd1 _06934_ sky130_fd_sc_hd__o22a_1
XFILLER_0_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_119_Left_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18265__Q team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[19\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16453_ clknet_leaf_180_wb_clk_i _02083_ _00149_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13665_ net2639 net240 net386 vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10877_ _06795_ _06873_ vssd1 vssd1 vccd1 vccd1 _06874_ sky130_fd_sc_hd__nor2_1
XANTENNA__09610__C net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12616_ _03651_ net1818 net202 vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__mux2_1
X_15404_ net1117 vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_119_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09075__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16384_ clknet_leaf_132_wb_clk_i _02014_ _00080_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13596_ net2261 net218 net395 vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18123_ clknet_leaf_47_wb_clk_i _00037_ _01819_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_15335_ net1199 vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__inv_2
X_12547_ _03662_ net1823 net205 vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__mux2_1
XANTENNA__12744__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08822__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18054_ net1039 _03392_ _01750_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_15266_ net1226 vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__inv_2
X_12478_ net1866 _03662_ net211 vssd1 vssd1 vccd1 vccd1 _03158_ sky130_fd_sc_hd__mux2_1
XANTENNA__10772__B _06768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_3 _06518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14217_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[13\] _04013_
+ _04014_ vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__o21a_1
X_17005_ clknet_leaf_159_wb_clk_i _02635_ _00701_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11429_ _07315_ _07319_ net1599 vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__o21ai_1
X_15197_ net1089 vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14148_ net1609 net506 net912 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[31\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_158_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13575__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15356__A net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14079_ _03925_ _03927_ _03945_ _03858_ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__a31o_1
X_17907_ clknet_leaf_75_wb_clk_i _03250_ _01603_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08889__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08353__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1070 net1071 vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__buf_4
Xfanout1081 net1086 vssd1 vssd1 vccd1 vccd1 net1081 sky130_fd_sc_hd__buf_4
X_08640_ _04710_ _04711_ _04712_ _04714_ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__or4_1
XFILLER_0_174_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17838_ clknet_leaf_78_wb_clk_i _03181_ _01534_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[84\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1092 net1094 vssd1 vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__buf_4
XFILLER_0_156_1060 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08571_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[25\]
+ net646 net619 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__a22o_1
X_17769_ clknet_leaf_99_wb_clk_i _03112_ _01465_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12919__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10999__A1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09123_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[12\]
+ net845 net785 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[12\]
+ _05178_ vssd1 vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08813__B1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout317_A _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08704__Y _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09054_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[13\]
+ net700 net597 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[13\]
+ _05112_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__a221o_1
XANTENNA__08433__A _04490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11130__Y _07096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold520 team_05_WB.instance_to_wrap.lcd_rs vssd1 vssd1 vccd1 vccd1 net1934 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_92_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold531 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 net1945 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap250 _03542_ vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_124_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1226_A net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold542 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 net1956 sky130_fd_sc_hd__dlygate4sd3_1
Xhold553 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[104\] vssd1 vssd1
+ vccd1 vccd1 net1967 sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[2\] vssd1 vssd1
+ vccd1 vccd1 net1978 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold575 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net1989 sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[10\] vssd1 vssd1
+ vccd1 vccd1 net2000 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08136__D_N team_05_WB.instance_to_wrap.total_design.data_from_keypad\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13485__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold597 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net2011 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08592__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09956_ net378 _04755_ vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_70_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1014_X net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08907_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[16\]
+ net687 net656 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__a22o_1
X_09887_ _04554_ _05915_ vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__nand2_4
XANTENNA_fanout474_X net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1220 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net2634 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout853_A _04367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1231 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2645 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1242 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2656 sky130_fd_sc_hd__dlygate4sd3_1
X_08838_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[18\]
+ net806 net760 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_142_Right_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1253 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2667 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1264 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net2678 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1275 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 net2689 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12428__A1 _07797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1286 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2700 sky130_fd_sc_hd__dlygate4sd3_1
X_08769_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[19\]
+ net676 net671 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout641_X net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1297 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2711 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12829__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout739_X net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10800_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[20\] team_05_WB.instance_to_wrap.total_design.core.program_count.imm_val_reg\[20\]
+ vssd1 vssd1 vccd1 vccd1 _06797_ sky130_fd_sc_hd__nand2_1
XANTENNA__10439__B1 _06280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_3__f_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09711__B net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11780_ _07573_ _07577_ _07578_ vssd1 vssd1 vccd1 vccd1 _07592_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09844__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18085__Q team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10731_ _06451_ net347 vssd1 vssd1 vccd1 vccd1 _06731_ sky130_fd_sc_hd__or2_1
XFILLER_0_165_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout906_X net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11651__A2 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_194_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_194_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_126_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13450_ net2124 net301 net415 vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__mux2_1
X_10662_ _05464_ net552 _06055_ _05812_ _06665_ vssd1 vssd1 vccd1 vccd1 _06666_ sky130_fd_sc_hd__o221a_1
XFILLER_0_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12401_ net1651 _07836_ _07852_ vssd1 vssd1 vccd1 vccd1 _03227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_123_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_123_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_91_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12600__A1 _07798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12564__S net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13381_ net2382 net278 net420 vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__mux2_1
X_10593_ _06593_ _06598_ _06600_ net536 vssd1 vssd1 vccd1 vccd1 _06601_ sky130_fd_sc_hd__a31o_1
XFILLER_0_118_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15120_ net1183 vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__inv_2
XANTENNA__10611__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12332_ net354 _03600_ _03626_ _03616_ _07510_ vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_114_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15051_ net1076 vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__inv_2
X_12263_ _07969_ _03557_ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14002_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[13\] _03847_ _03845_
+ vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__a21o_1
X_11214_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[13\] _07101_
+ _07127_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[125\] vssd1
+ vssd1 vccd1 vccd1 _07178_ sky130_fd_sc_hd__a22o_1
X_12194_ _08005_ _07982_ _07983_ vssd1 vssd1 vccd1 vccd1 _08006_ sky130_fd_sc_hd__mux2_2
XANTENNA__13395__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15176__A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08583__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11145_ _07038_ _07075_ _07079_ vssd1 vssd1 vccd1 vccd1 _07111_ sky130_fd_sc_hd__and3_4
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__clkbuf_4
X_11076_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[4\] team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[3\]
+ vssd1 vssd1 vccd1 vccd1 _07043_ sky130_fd_sc_hd__or2_1
X_15953_ net1269 vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__inv_2
XANTENNA__09605__C net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12312__B _03605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10027_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[13\] _06055_
+ vssd1 vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__nor2_2
X_14904_ net1210 vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__inv_2
X_15884_ net1293 vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__inv_2
X_17623_ clknet_leaf_59_wb_clk_i _02994_ _01319_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_14835_ net1213 vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__inv_2
XANTENNA__12739__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_127_Left_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09180__Y _05234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17554_ clknet_leaf_65_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[25\]
+ _01250_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11978_ net501 _07684_ vssd1 vssd1 vccd1 vccd1 _07790_ sky130_fd_sc_hd__nor2_1
X_14766_ net1180 vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09296__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10767__B _06764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09835__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16505_ clknet_leaf_15_wb_clk_i _02135_ _00201_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13717_ net905 _06464_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[17\]
+ sky130_fd_sc_hd__and2_1
X_10929_ _06878_ _06919_ vssd1 vssd1 vccd1 vccd1 _06920_ sky130_fd_sc_hd__xnor2_1
X_17485_ clknet_leaf_36_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[20\]
+ _01181_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_14697_ net1215 vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__inv_2
XFILLER_0_160_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08237__B net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09048__B1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16436_ clknet_leaf_120_wb_clk_i _02066_ _00132_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13648_ net2593 net298 net390 vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11879__A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09599__A1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13579_ net2090 net278 net396 vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__mux2_1
X_16367_ clknet_leaf_135_wb_clk_i _01997_ _00063_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13797__C net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18106_ clknet_leaf_55_wb_clk_i _03429_ _01802_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_15318_ net1084 vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__inv_2
X_16298_ net1148 vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_136_Left_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18037_ clknet_leaf_94_wb_clk_i _03375_ _01733_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_10_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15249_ net1192 vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09636__X team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09220__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09810_ _04879_ _05840_ _04881_ vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__a21oi_4
Xfanout307 net308 vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__buf_2
XANTENNA__08574__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout318 _06671_ vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__buf_1
Xfanout329 _06705_ vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__dlymetal6s2s_1
X_09741_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[0\]
+ net880 net873 net866 vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__and4_1
XFILLER_0_158_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09672_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[1\]
+ net876 net860 net857 vssd1 vssd1 vccd1 vccd1 _05705_ sky130_fd_sc_hd__and4_1
XFILLER_0_94_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_145_Left_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08623_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[24\]
+ net834 net749 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08554_ _04616_ _04617_ _04629_ _04630_ vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__or4_1
XANTENNA__09287__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09826__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11125__Y _07091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11633__A2 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08485_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[27\]
+ net713 net684 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[27\]
+ _04562_ vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout434_A _03722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1176_A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09039__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12384__S _03660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12594__A0 _03632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09106_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[12\]
+ net699 net644 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[12\]
+ _05147_ vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09037_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[14\]
+ net848 _05094_ _05096_ net856 vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__a2111o_1
XANTENNA__14335__B2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold350 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[38\] vssd1 vssd1
+ vccd1 vccd1 net1764 sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[80\] vssd1 vssd1
+ vccd1 vccd1 net1775 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09211__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout591_X net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold372 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[82\] vssd1 vssd1
+ vccd1 vccd1 net1786 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout689_X net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold383 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[60\] vssd1 vssd1
+ vccd1 vccd1 net1797 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08565__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold394 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1808 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout830 net832 vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__clkbuf_8
Xfanout841 net844 vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__clkbuf_8
Xfanout852 _04370_ vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__buf_2
X_09939_ _05035_ _05055_ _05967_ vssd1 vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout856_X net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout863 _04294_ vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__buf_2
Xfanout874 net875 vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__buf_2
XANTENNA__11029__A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout885 _04281_ vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__clkbuf_2
Xfanout896 net898 vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__clkbuf_2
X_12950_ net290 net2502 net468 vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__mux2_1
Xhold1050 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 net2464 sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ _07710_ _07712_ vssd1 vssd1 vccd1 vccd1 _07713_ sky130_fd_sc_hd__and2_1
Xhold1061 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1072 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net2486 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12881_ net280 net2501 net476 vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__mux2_1
Xhold1083 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2497 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12559__S net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1094 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 net2508 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14620_ net1083 vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11832_ _07633_ _07634_ _07642_ _07643_ _07619_ vssd1 vssd1 vccd1 vccd1 _07644_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_169_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09817__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14551_ net1104 vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__inv_2
X_11763_ _07547_ _07560_ _07574_ vssd1 vssd1 vccd1 vccd1 _07575_ sky130_fd_sc_hd__o21a_1
XANTENNA__10079__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13502_ net2389 net230 net405 vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__mux2_1
X_10714_ net332 _06582_ _06712_ net335 _06714_ vssd1 vssd1 vccd1 vccd1 _06715_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_155_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17270_ clknet_leaf_139_wb_clk_i _02900_ _00966_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14482_ net1239 vssd1 vssd1 vccd1 vccd1 _00112_ sky130_fd_sc_hd__inv_2
X_11694_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[27\] net1000 vssd1
+ vssd1 vccd1 vccd1 _07506_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16221_ net1054 vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__inv_2
X_13433_ net1947 net243 net415 vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__mux2_1
X_10645_ net332 _06506_ net347 _06360_ _06648_ vssd1 vssd1 vccd1 vccd1 _06650_ sky130_fd_sc_hd__o221a_1
XANTENNA__12585__A0 _03657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16152_ net1153 vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13364_ net2021 net191 net422 vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__mux2_1
X_10576_ _06576_ _06583_ _06584_ net536 vssd1 vssd1 vccd1 vccd1 _06585_ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09450__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12315_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[21\] net1000 _08022_
+ _03609_ net544 vssd1 vssd1 vccd1 vccd1 _03610_ sky130_fd_sc_hd__a221o_4
XANTENNA__11986__X _07798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15103_ net1182 vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__inv_2
X_16083_ net1259 vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__inv_2
XANTENNA__14326__B2 _05165_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13295_ _04252_ _04254_ _04255_ _04259_ vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__and4_1
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10108__A _05165_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1032 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15034_ net1058 vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__inv_2
X_12246_ _03536_ _03540_ vssd1 vssd1 vccd1 vccd1 _03541_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_91_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_82_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08556__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[26\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12352__A3 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[12\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12177_ _07933_ _07937_ _07939_ _07931_ vssd1 vssd1 vccd1 vccd1 _07989_ sky130_fd_sc_hd__or4b_1
XANTENNA__09616__B net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_20_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11128_ _07093_ vssd1 vssd1 vccd1 vccd1 _07094_ sky130_fd_sc_hd__inv_2
X_16985_ clknet_leaf_5_wb_clk_i _02615_ _00681_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11059_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[1\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[0\]
+ vssd1 vssd1 vccd1 vccd1 _07026_ sky130_fd_sc_hd__nand2_1
X_15936_ net1265 vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12469__S net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15867_ net1304 vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17606_ clknet_leaf_81_wb_clk_i _02977_ _01302_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14818_ net1216 vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09269__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15798_ net1297 vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__inv_2
XANTENNA__10497__B net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17537_ clknet_leaf_81_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[8\]
+ _01233_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11615__A2 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14749_ net1089 vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08270_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[30\] team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[20\]
+ _04352_ vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__nor3_2
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17468_ clknet_leaf_41_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[3\]
+ _01164_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_2__f_wb_clk_i_X clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16419_ clknet_leaf_199_wb_clk_i _02049_ _00115_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17399_ clknet_leaf_59_wb_clk_i net1431 _01095_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg2\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12576__A0 _03623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14317__A1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08795__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12932__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14317__B2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[18\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08547__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10354__A2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout384_A net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09724_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[0\]
+ net768 _05748_ _05751_ _05753_ vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__a2111oi_1
XTAP_TAPCELL_ROW_87_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09655_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[1\]
+ net846 net841 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[1\]
+ _05680_ vssd1 vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__a221o_1
XANTENNA__12379__S net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10688__A net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout551_A net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11136__X _07102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout649_A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08606_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[24\]
+ net689 net681 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_26_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09586_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[2\]
+ net1015 net943 net927 vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__and4_1
XFILLER_0_171_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08537_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[26\]
+ net835 net828 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout816_A _04388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout437_X net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08468_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[28\]
+ net789 net758 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08399_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[29\]
+ net607 net597 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[29\]
+ _04478_ vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout604_X net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13003__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10430_ net892 _06445_ _06444_ _05924_ vssd1 vssd1 vccd1 vccd1 _06446_ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09432__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12127__B _07657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08324__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10361_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[21\] _06097_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06381_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12842__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12100_ _07902_ _07910_ _07864_ vssd1 vssd1 vccd1 vccd1 _07912_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13080_ net282 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[13\]
+ net452 vssd1 vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__mux2_1
X_10292_ net895 _06314_ vssd1 vssd1 vccd1 vccd1 _06315_ sky130_fd_sc_hd__nor2_1
XANTENNA__14342__B team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12031_ _07450_ _07842_ vssd1 vssd1 vccd1 vccd1 _07843_ sky130_fd_sc_hd__nor2_2
XANTENNA__08538__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold180 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i_reg\[23\]
+ vssd1 vssd1 vccd1 vccd1 net1594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[15\] vssd1 vssd1
+ vccd1 vccd1 net1605 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08340__B net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout660 net663 vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11982__A _07789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13673__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout671 _04304_ vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__clkbuf_8
X_16770_ clknet_leaf_7_wb_clk_i _02400_ _00466_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout682 _04301_ vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__clkbuf_8
X_13982_ _03852_ _03853_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__nand2b_1
XANTENNA__09499__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout693 net694 vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__buf_4
X_15721_ net1142 vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_126_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12933_ net220 net2531 net470 vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_126_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10598__A net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08710__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15652_ net1243 vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12864_ net190 net2539 net478 vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__mux2_1
XANTENNA__09602__D net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14603_ net1067 vssd1 vssd1 vccd1 vccd1 _00233_ sky130_fd_sc_hd__inv_2
X_18371_ net1356 vssd1 vssd1 vccd1 vccd1 la_data_out[19] sky130_fd_sc_hd__buf_2
X_11815_ _07607_ _07626_ vssd1 vssd1 vccd1 vccd1 _07627_ sky130_fd_sc_hd__and2_2
X_15583_ net1251 vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12795_ _04261_ net562 _03702_ vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__or3_4
XFILLER_0_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13702__A net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17322_ clknet_leaf_181_wb_clk_i _02952_ _01018_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11746_ _07554_ _07555_ _07557_ vssd1 vssd1 vccd1 vccd1 _07558_ sky130_fd_sc_hd__a21o_1
X_14534_ net1231 vssd1 vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_174_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_174_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18273__Q team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[27\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17253_ clknet_leaf_180_wb_clk_i _02883_ _00949_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11677_ _07491_ vssd1 vssd1 vccd1 vccd1 _07492_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_12_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14465_ net1235 vssd1 vssd1 vccd1 vccd1 _00095_ sky130_fd_sc_hd__inv_2
XANTENNA__12558__A0 _03614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16204_ net1079 vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10628_ _06625_ _06626_ _06633_ net537 vssd1 vssd1 vccd1 vccd1 _06634_ sky130_fd_sc_hd__a31o_1
X_13416_ net2146 net288 net416 vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14396_ net1488 vssd1 vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17184_ clknet_leaf_132_wb_clk_i _02814_ _00880_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09423__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08234__C _04287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11230__B1 _07169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16135_ net1310 vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08777__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13347_ net282 net2283 net425 vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__mux2_1
X_10559_ net898 _06568_ vssd1 vssd1 vccd1 vccd1 _06569_ sky130_fd_sc_hd__nor2_1
XANTENNA__12752__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_51_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10584__A2 _06591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16066_ net1173 vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__inv_2
X_13278_ net268 net2629 net432 vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08529__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12229_ _03521_ _03522_ _03518_ _03519_ vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__a2bb2o_2
X_15017_ net1222 vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__inv_2
XANTENNA__10272__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13583__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16968_ clknet_leaf_197_wb_clk_i _02598_ _00664_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11297__B1 _07113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15919_ net1302 vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10639__A3 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16899_ clknet_leaf_199_wb_clk_i _02529_ _00595_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08701__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09440_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[5\]
+ net718 _05479_ _05482_ vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_148_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09371_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[7\]
+ net819 net807 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[7\]
+ _05401_ vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_82_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08322_ net942 net935 net932 vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_58_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_74_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09662__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08253_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[31\]
+ net634 net603 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__a22o_1
XANTENNA__10447__S net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14146__C net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08184_ _04233_ net958 vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__nand2_2
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09414__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10024__A1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11221__B1 _07119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10575__A2 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17527__Q team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[30\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout599_A net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1306_A net1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09193__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout387_X net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout766_A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08940__A2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11288__B1 _07130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09707_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[24\]\[0\]
+ net950 net939 net936 vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__and4_1
XANTENNA_clkbuf_leaf_97_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout933_A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout554_X net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09638_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[1\]
+ net946 net930 net924 vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__and4_1
XFILLER_0_167_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08319__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout721_X net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09569_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[2\]
+ net941 net1013 net932 vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__and4_1
XANTENNA__12837__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout819_X net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11600_ net1644 net1009 net345 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12580_ _03661_ net1816 net203 vssd1 vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09653__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11531_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write
+ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[13\] vssd1 vssd1 vccd1
+ vccd1 _07442_ sky130_fd_sc_hd__o21a_1
XFILLER_0_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08335__B net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14250_ team_05_WB.instance_to_wrap.total_design.keypad0.counter\[7\] _04020_ vssd1
+ vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11462_ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[7\] _07372_ net1002
+ vssd1 vssd1 vccd1 vccd1 _07373_ sky130_fd_sc_hd__mux2_2
XFILLER_0_135_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09405__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13201_ net235 net2246 net352 vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__mux2_1
XANTENNA__11212__B1 _07169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08759__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire379 _04697_ vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13668__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10413_ _06395_ _06429_ net519 vssd1 vssd1 vccd1 vccd1 _06430_ sky130_fd_sc_hd__mux2_1
X_14181_ net1923 net503 net908 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[30\]
+ sky130_fd_sc_hd__and3_1
X_11393_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[7\] team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_20ms\[6\]
+ _07323_ vssd1 vssd1 vccd1 vccd1 _07324_ sky130_fd_sc_hd__and3_1
XANTENNA__12572__S _03678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_204_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_61_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13132_ net223 net2742 net445 vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input62_A wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10344_ team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[23\] net903 net965
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 _06365_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_78_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17940_ clknet_leaf_34_wb_clk_i _03279_ _01636_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13063_ net196 net2171 net454 vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__mux2_1
X_10275_ net525 _06205_ vssd1 vssd1 vccd1 vccd1 _06298_ sky130_fd_sc_hd__or2_1
X_12014_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[31\] team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[23\]
+ net995 net548 vssd1 vssd1 vccd1 vccd1 _07826_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_167_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17871_ clknet_leaf_89_wb_clk_i _03214_ _01567_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_output149_A net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08392__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08931__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16822_ clknet_leaf_151_wb_clk_i _02452_ _00518_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout490 _03700_ vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11279__B1 _07121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18268__Q team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[22\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16753_ clknet_leaf_118_wb_clk_i _02383_ _00449_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13965_ net2972 net507 _03837_ vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__a21oi_1
X_15704_ net1166 vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__inv_2
X_12916_ net289 net2673 net472 vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__mux2_1
X_16684_ clknet_leaf_7_wb_clk_i _02314_ _00380_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10121__A _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13896_ net1559 net981 _03784_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[19\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_100_Left_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09910__A _05350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15635_ net1245 vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__inv_2
XANTENNA__12747__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12847_ net284 net2703 net482 vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__mux2_1
XANTENNA__12779__A0 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18354_ net1339 vssd1 vssd1 vccd1 vccd1 la_data_out[2] sky130_fd_sc_hd__buf_2
X_15566_ net1244 vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12778_ net275 net2341 net491 vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17305_ clknet_leaf_15_wb_clk_i _02935_ _01001_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14517_ net1059 vssd1 vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11729_ team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[10\] net997 vssd1
+ vssd1 vccd1 vccd1 _07541_ sky130_fd_sc_hd__nand2_1
X_18285_ net1377 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
XFILLER_0_16_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15497_ net1156 vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17236_ clknet_leaf_112_wb_clk_i _02866_ _00932_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14448_ net1195 vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13578__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12482__S net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17167_ clknet_leaf_139_wb_clk_i _02797_ _00863_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14379_ net1501 vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold905 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 net2319 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold916 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[5\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 net2330 sky130_fd_sc_hd__dlygate4sd3_1
Xhold927 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2341 sky130_fd_sc_hd__dlygate4sd3_1
X_16118_ net1134 vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__inv_2
Xhold938 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net2352 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08261__A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold949 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2363 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17098_ clknet_leaf_17_wb_clk_i _02728_ _00794_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08940_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[16\]
+ net841 net786 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__a22o_1
X_16049_ net1285 vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__inv_2
XANTENNA__09175__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_131_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08871_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[17\]
+ net628 net607 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[17\]
+ _04937_ vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__a221o_1
XANTENNA__10015__B net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08922__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09423_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[5\]
+ net702 net639 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14438__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09354_ _05400_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[7\]
+ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1089_A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09635__B1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[21\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10685__B _06687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10245__A1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[27\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08305_ net945 net1013 net933 vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__and3_1
XANTENNA__11133__Y _07099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08989__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09285_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[8\]
+ net650 net623 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[8\]
+ _05333_ vssd1 vssd1 vccd1 vccd1 _05334_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout514_A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08236_ net883 net871 net864 vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__and3_4
XFILLER_0_7_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13488__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12392__S _07852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08167_ team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[8\] _04249_
+ vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_170_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_31_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08098_ net1036 net1019 net975 _04198_ vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_56_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08171__A team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[10\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout883_A net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1211_X net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09166__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_148_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_148_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10060_ team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[8\] _06088_ vssd1
+ vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_73_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_73_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout671_X net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17634__D team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08374__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout769_X net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08913__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09714__B net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout936_X net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09323__C1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13750_ _05212_ _06445_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[18\]
+ sky130_fd_sc_hd__and2_1
X_10962_ _06439_ _06768_ net564 vssd1 vssd1 vccd1 vccd1 _06947_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12701_ net231 net2419 net497 vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__mux2_1
XANTENNA__12567__S _03678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10893_ net1044 _06104_ net957 vssd1 vssd1 vccd1 vccd1 _06890_ sky130_fd_sc_hd__o21a_1
X_13681_ net2329 net300 net385 vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__mux2_1
XANTENNA__11471__S net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15420_ net1124 vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__inv_2
X_12632_ _03664_ net1907 net202 vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08346__A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12563_ net1752 _03663_ _03678_ vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15351_ net1103 vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11514_ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[23\] _07424_ net1003
+ vssd1 vssd1 vccd1 vccd1 _07425_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14302_ _04533_ _04552_ vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__and2_1
X_18070_ clknet_leaf_85_wb_clk_i _00006_ _01766_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12494_ net1734 _03663_ _03673_ vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15282_ net1238 vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13398__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17021_ clknet_leaf_110_wb_clk_i _02651_ _00717_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11445_ team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[30\] _07356_ net1003
+ vssd1 vssd1 vccd1 vccd1 _07357_ sky130_fd_sc_hd__mux2_1
X_14233_ team_05_WB.instance_to_wrap.total_design.keypad0.counter\[16\] _04026_ net2323
+ vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_169_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14164_ _03992_ net907 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[13\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_169_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11376_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[4\] _07072_
+ net731 vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09608__C net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_156_Right_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10327_ _05983_ _05986_ _05929_ vssd1 vssd1 vccd1 vccd1 _06348_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13115_ net290 net2804 net448 vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__mux2_1
X_14095_ _03961_ _03858_ _03960_ vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__or3b_1
XANTENNA__14811__A net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17923_ clknet_leaf_43_wb_clk_i _03262_ _01619_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.CPU_DAT_O\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13046_ net276 net2858 net458 vssd1 vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__mux2_1
XANTENNA__09905__A _04989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10258_ _06164_ _06174_ vssd1 vssd1 vccd1 vccd1 _06282_ sky130_fd_sc_hd__nand2_1
Xfanout1230 net1234 vssd1 vssd1 vccd1 vccd1 net1230 sky130_fd_sc_hd__buf_4
Xfanout1241 net1313 vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__buf_4
X_17854_ clknet_leaf_76_wb_clk_i _03197_ _01550_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[36\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1252 net1312 vssd1 vssd1 vccd1 vccd1 net1252 sky130_fd_sc_hd__buf_2
X_10189_ net897 _06214_ _06215_ _06213_ vssd1 vssd1 vccd1 vccd1 _06216_ sky130_fd_sc_hd__o211ai_2
Xfanout1263 net1264 vssd1 vssd1 vccd1 vccd1 net1263 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1274 net1278 vssd1 vssd1 vccd1 vccd1 net1274 sky130_fd_sc_hd__clkbuf_2
X_16805_ clknet_leaf_22_wb_clk_i _02435_ _00501_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1285 net1286 vssd1 vssd1 vccd1 vccd1 net1285 sky130_fd_sc_hd__buf_2
Xfanout1296 net1298 vssd1 vssd1 vccd1 vccd1 net1296 sky130_fd_sc_hd__buf_2
X_17785_ clknet_leaf_99_wb_clk_i _03128_ _01481_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_14997_ net1060 vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__inv_2
XFILLER_0_163_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16736_ clknet_leaf_132_wb_clk_i _02366_ _00432_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[18\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13948_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[6\] team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__nand2_1
XANTENNA__08808__X team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[19\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12477__S net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16667_ clknet_leaf_190_wb_clk_i _02297_ _00363_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13879_ team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_reg\[11\]
+ net561 net575 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_reg\[11\]
+ net986 vssd1 vssd1 vccd1 vccd1 _03776_ sky130_fd_sc_hd__a221o_1
X_18406_ net914 vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15618_ net1157 vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__inv_2
XANTENNA__13413__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16598_ clknet_leaf_142_wb_clk_i _02228_ _00294_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18337_ net1326 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
XFILLER_0_17_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15549_ net1124 vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09070_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[6\]\[13\]
+ net832 net795 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18268_ clknet_leaf_33_wb_clk_i _03497_ _01963_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_47_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17219_ clknet_leaf_196_wb_clk_i _02849_ _00915_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18199_ clknet_leaf_33_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_out_INSTR\[20\]
+ _01894_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_i\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12924__A0 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold702 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[2\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2116 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13101__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold713 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 net2127 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold724 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 net2138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2160 sky130_fd_sc_hd__dlygate4sd3_1
Xhold757 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 net2182 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10026__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09972_ net891 _06000_ _05924_ _05922_ vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__o211a_1
XANTENNA__12940__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold779 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 net2193 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09148__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08923_ _04973_ _04974_ _04986_ _04987_ vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__or4_1
XANTENNA__08356__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_51_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1402 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net2816 sky130_fd_sc_hd__dlygate4sd3_1
X_08854_ net571 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[18\]
+ team_05_WB.instance_to_wrap.total_design.core.ctrl.imm_32\[18\] vssd1 vssd1 vccd1
+ vccd1 _04921_ sky130_fd_sc_hd__a21oi_1
Xhold1413 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 net2827 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1424 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 net2838 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1435 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net2849 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1446 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[3\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 net2860 sky130_fd_sc_hd__dlygate4sd3_1
X_08785_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[7\]\[19\]
+ net660 _04855_ net719 vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__a211o_1
XFILLER_0_58_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1457 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 net2871 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1468 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[14\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1479 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2893 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout464_A _03710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10466__A1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09320__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12387__S _07852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout631_A _04314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout729_A net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09406_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[6\]
+ net799 net765 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[22\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09337_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[12\]\[7\]
+ net696 net677 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1161_X net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09268_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[9\]
+ net803 net799 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05318_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08219_ net878 net869 net858 vssd1 vssd1 vccd1 vccd1 _04302_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09709__B net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09199_ _05245_ _05247_ _05249_ _05251_ vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__or4_1
XFILLER_0_133_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13011__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11230_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[100\] _07123_
+ _07169_ _07192_ vssd1 vssd1 vccd1 vccd1 _07193_ sky130_fd_sc_hd__a211o_1
XFILLER_0_160_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09387__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12391__A1 _07798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11194__A2 _07104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11161_ _07039_ _07098_ vssd1 vssd1 vccd1 vccd1 _07127_ sky130_fd_sc_hd__nor2_4
XFILLER_0_31_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12850__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10941__A2 _06768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18364__1349 vssd1 vssd1 vccd1 vccd1 _18364__1349/HI net1349 sky130_fd_sc_hd__conb_1
XANTENNA__09139__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10112_ _06132_ _06139_ net528 vssd1 vssd1 vccd1 vccd1 _06140_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11092_ _07052_ _07058_ vssd1 vssd1 vccd1 vccd1 _07059_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_164_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14920_ net1223 vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__inv_2
X_10043_ net521 _06069_ _06071_ _06060_ net531 vssd1 vssd1 vccd1 vccd1 _06072_ sky130_fd_sc_hd__o2111a_1
XANTENNA__10154__B1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold40 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[13\]
+ vssd1 vssd1 vccd1 vccd1 net1454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[9\]
+ vssd1 vssd1 vccd1 vccd1 net1465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[31\] vssd1 vssd1
+ vccd1 vccd1 net1476 sky130_fd_sc_hd__dlygate4sd3_1
X_14851_ net1200 vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__inv_2
XANTENNA_input25_A DAT_I[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold73 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[10\]
+ vssd1 vssd1 vccd1 vccd1 net1487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[14\] vssd1 vssd1
+ vccd1 vccd1 net1498 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13681__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold95 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[6\]
+ vssd1 vssd1 vccd1 vccd1 net1509 sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ net1567 net977 net725 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[13\]
+ sky130_fd_sc_hd__and3_1
X_17570_ clknet_leaf_114_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[7\]
+ _01266_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14782_ net1054 vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__inv_2
X_11994_ net356 _07565_ _07768_ _07796_ vssd1 vssd1 vccd1 vccd1 _07806_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_98_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09311__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16521_ clknet_leaf_20_wb_clk_i _02151_ _00217_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13733_ net922 _06743_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_write_adr_i\[1\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__10457__B2 _06355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10945_ net1042 _06382_ net956 vssd1 vssd1 vccd1 vccd1 _06933_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_45_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_156_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16452_ clknet_leaf_194_wb_clk_i _02082_ _00148_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[27\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13664_ net1983 net243 net386 vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__mux2_1
X_10876_ _06798_ _06872_ _06797_ vssd1 vssd1 vccd1 vccd1 _06873_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_73_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09610__D net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15403_ net1138 vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12615_ _03662_ net1898 net202 vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__mux2_1
XANTENNA__13946__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16383_ clknet_leaf_156_wb_clk_i _02013_ _00079_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[29\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13595_ net2267 net189 net393 vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18122_ clknet_leaf_47_wb_clk_i _00036_ _01818_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15334_ net1230 vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__inv_2
X_12546_ _03661_ net1938 net205 vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18053_ net1039 _03391_ _01749_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_15265_ net1225 vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__inv_2
XANTENNA__10545__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12477_ net1744 _03661_ net210 vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_4 _06518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17004_ clknet_leaf_2_wb_clk_i _02634_ _00700_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_14216_ team_05_WB.instance_to_wrap.total_design.lcd_display.cnt_500hz\[13\] _04013_
+ net728 vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__a21boi_1
X_11428_ _07313_ _07342_ net730 vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__a21o_1
X_15196_ net1064 vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__inv_2
XANTENNA__11185__A2 _07115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12382__A1 _03612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08586__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11359_ _07300_ team_05_WB.instance_to_wrap.total_design.keypad0.key_out\[2\] net509
+ vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__mux2_1
X_14147_ net1923 net503 net911 vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_bus_i\[30\]
+ sky130_fd_sc_hd__and3_1
X_14078_ _03925_ _03927_ _03945_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08338__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11376__S net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17906_ clknet_leaf_91_wb_clk_i _03249_ _01602_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13029_ net200 net2909 net459 vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__mux2_1
Xfanout1060 net1061 vssd1 vssd1 vccd1 vccd1 net1060 sky130_fd_sc_hd__buf_4
Xfanout1071 net1072 vssd1 vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__buf_4
X_17837_ clknet_leaf_101_wb_clk_i _03180_ _01533_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[83\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09550__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1082 net1086 vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__clkbuf_4
Xfanout1093 net1094 vssd1 vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13591__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15372__A net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08570_ _04639_ _04641_ _04643_ _04645_ vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__or4_1
XFILLER_0_156_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17768_ clknet_leaf_90_wb_clk_i _03111_ _01464_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16719_ clknet_leaf_135_wb_clk_i _02349_ _00415_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_17699_ clknet_leaf_89_wb_clk_i _03042_ _01395_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.lcd_display.row_1\[73\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08510__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11124__B net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12935__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09122_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[12\]
+ net826 net825 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_44_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09053_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[15\]\[13\]
+ net665 net640 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[11\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_96_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout212_A net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09369__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold510 net104 vssd1 vssd1 vccd1 vccd1 net1924 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold521 net106 vssd1 vssd1 vccd1 vccd1 net1935 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10027__Y _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12373__A1 _07791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11176__A2 _07108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08577__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold532 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[26\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1946 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap251 _03550_ vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__clkbuf_2
Xhold543 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 net1957 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold554 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[21\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 net1968 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold565 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[13\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1979 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1121_A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold576 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 net1990 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold587 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[23\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2001 sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 team_05_WB.instance_to_wrap.total_design.core.data_bus_o\[8\] vssd1 vssd1
+ vccd1 vccd1 net2012 sky130_fd_sc_hd__dlygate4sd3_1
X_09955_ _05977_ _05978_ _05979_ _05982_ _05929_ vssd1 vssd1 vccd1 vccd1 _05984_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_70_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout581_A net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08906_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[16\]
+ net652 net636 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__a22o_1
X_09886_ _04533_ _04553_ vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__or2_1
Xhold1210 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 net2624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1221 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[10\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 net2635 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09541__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1232 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[1\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2646 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08837_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[18\]
+ net833 net826 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[31\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__a22o_1
Xhold1243 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[8\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 net2657 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1254 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[16\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 net2668 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout846_A _04373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout467_X net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1265 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[17\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 net2679 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1276 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 net2690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1287 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[4\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 net2701 sky130_fd_sc_hd__dlygate4sd3_1
X_08768_ _04818_ _04838_ vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__nand2_1
Xhold1298 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[9\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 net2712 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10439__A1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10439__B2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout634_X net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09711__C net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08699_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[20\]\[22\]
+ net599 _04771_ net721 vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__a211o_1
XANTENNA__13006__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10730_ net888 _06729_ _06728_ vssd1 vssd1 vccd1 vccd1 _06730_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10661_ net524 _06663_ _06664_ vssd1 vssd1 vccd1 vccd1 _06665_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_24_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12845__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout801_X net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12400_ net1672 _03650_ net217 vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__mux2_1
XANTENNA__11602__X _07474_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09279__X team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13380_ net2059 net283 net420 vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__mux2_1
X_10592_ _06049_ _06279_ _06597_ _06599_ vssd1 vssd1 vccd1 vccd1 _06600_ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12331_ net250 net251 _03591_ _03601_ vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_133_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_163_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_163_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12262_ _07951_ _03555_ _03556_ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__a21o_1
X_15050_ net1110 vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__inv_2
XANTENNA__11167__A2 _07105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11213_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[93\] _07096_
+ _07123_ team_05_WB.instance_to_wrap.total_design.lcd_display.row_2\[101\] _07176_
+ vssd1 vssd1 vccd1 vccd1 _07177_ sky130_fd_sc_hd__a221o_1
X_14001_ _03867_ _03870_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08568__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13676__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12580__S net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12193_ _07982_ _07985_ vssd1 vssd1 vccd1 vccd1 _08005_ sky130_fd_sc_hd__nand2_1
X_11144_ _07083_ _07087_ vssd1 vssd1 vccd1 vccd1 _07110_ sky130_fd_sc_hd__nor2_4
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__clkbuf_4
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__clkbuf_4
X_11075_ team_05_WB.instance_to_wrap.total_design.lcd_display.currentState\[3\] _07041_
+ vssd1 vssd1 vccd1 vccd1 _07042_ sky130_fd_sc_hd__nor2_1
X_15952_ net1266 vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__inv_2
XANTENNA__11324__C1 _07031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09605__D net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10026_ net1018 _05923_ vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__or2_2
X_14903_ net1096 vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__inv_2
XANTENNA__09532__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output131_A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15883_ net1303 vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__inv_2
XANTENNA__08740__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17622_ clknet_leaf_64_wb_clk_i _02993_ _01318_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.instr_mem.instruction_adr_stored\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13705__A net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14834_ net1240 vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17553_ clknet_leaf_63_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_data_adr\[24\]
+ _01249_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_adr_o\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__18276__Q team_05_WB.instance_to_wrap.total_design.core.ctrl.instruction\[30\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14765_ net1087 vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__inv_2
X_11977_ _07788_ _07787_ _07518_ _07506_ vssd1 vssd1 vccd1 vccd1 _07789_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_98_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16504_ clknet_leaf_29_wb_clk_i _02134_ _00200_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[25\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13716_ _04235_ _06481_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_read_adr_i\[16\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10928_ _06786_ _06787_ vssd1 vssd1 vccd1 vccd1 _06919_ sky130_fd_sc_hd__or2_1
X_17484_ clknet_leaf_36_wb_clk_i team_05_WB.instance_to_wrap.total_design.core.data_mem.stored_read_data\[19\]
+ _01180_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.data_cpu_o\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_14696_ net1218 vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08237__C net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10850__A1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16435_ clknet_leaf_164_wb_clk_i _02065_ _00131_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[28\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13919__A2 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12755__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13647_ net2174 net288 net388 vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__mux2_1
X_10859_ _06825_ _06855_ vssd1 vssd1 vccd1 vccd1 _06856_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14337__A2_N team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[15\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09599__A2 team_05_WB.instance_to_wrap.total_design.core.data_mem.data_cpu_i\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10666__A2_N net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11879__B _07690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16366_ clknet_leaf_171_wb_clk_i _01996_ _00062_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.regFile.register\[30\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13578_ net2244 net283 net396 vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__mux2_1
X_18105_ clknet_leaf_53_wb_clk_i _03428_ _01801_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.total_design.core.math.pc_val\[22\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_54_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15317_ net1059 vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__inv_2
X_12529_ net1697 _03664_ net209 vssd1 vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__mux2_1
X_16297_ net1148 vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18036_ clknet_leaf_43_wb_clk_i net1469 _01732_ vssd1 vssd1 vccd1 vccd1 team_05_WB.instance_to_wrap.wishbone.prev_BUSY_O
+ sky130_fd_sc_hd__dfrtp_1
X_15248_ net1093 vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13586__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12490__S net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15179_ net1071 vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout308 _06767_ vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__clkbuf_2
Xfanout319 _06671_ vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__buf_2
X_09740_ team_05_WB.instance_to_wrap.total_design.core.regFile.register\[19\]\[0\]
+ net886 net873 net868 vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__and4_1
.ends

