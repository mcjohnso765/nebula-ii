* NGSPICE file created from team_01_Wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_16 abstract view
.subckt sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_1 abstract view
.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_2 abstract view
.subckt sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

.subckt team_01_Wrapper ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14]
+ ADR_O[15] ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22]
+ ADR_O[23] ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30]
+ ADR_O[31] ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0]
+ DAT_I[10] DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17]
+ DAT_I[18] DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25]
+ DAT_I[26] DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4]
+ DAT_I[5] DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12]
+ DAT_O[13] DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20]
+ DAT_O[21] DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28]
+ DAT_O[29] DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7]
+ DAT_O[8] DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[34] gpio_in[35] gpio_in[36]
+ gpio_in[37] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9]
+ gpio_oeb[0] gpio_oeb[10] gpio_oeb[11] gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15]
+ gpio_oeb[16] gpio_oeb[17] gpio_oeb[18] gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21]
+ gpio_oeb[22] gpio_oeb[23] gpio_oeb[24] gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28]
+ gpio_oeb[29] gpio_oeb[2] gpio_oeb[30] gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[34]
+ gpio_oeb[35] gpio_oeb[36] gpio_oeb[37] gpio_oeb[3] gpio_oeb[4] gpio_oeb[5] gpio_oeb[6]
+ gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12]
+ gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19]
+ gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25]
+ gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31]
+ gpio_out[32] gpio_out[33] gpio_out[34] gpio_out[35] gpio_out[36] gpio_out[37] gpio_out[3]
+ gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] irq[0] irq[1]
+ irq[2] la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13]
+ la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19]
+ la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24]
+ la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2]
+ la_data_in[30] la_data_in[31] la_data_in[3] la_data_in[4] la_data_in[5] la_data_in[6]
+ la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10] la_data_out[11]
+ la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16]
+ la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21]
+ la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26]
+ la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31]
+ la_data_out[3] la_data_out[4] la_data_out[5] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[3] la_oenb[4]
+ la_oenb[5] la_oenb[6] la_oenb[7] la_oenb[8] la_oenb[9] vccd1 vssd1 wb_clk_i wb_rst_i
+ wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XANTENNA__09523__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09671_ net993 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[22\] _04662_
+ vssd1 vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11834__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08622_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[11\] net662 net658 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__a22o_1
XANTENNA__13607__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08709__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11618__A0 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08553_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[19\] net661 _04890_
+ _04891_ _04892_ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_77_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09531__C net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08428__B net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08484_ net1081 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[23\] net887
+ vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__and3_1
XANTENNA__14017__D1 _04152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10841__A1 _06098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12665__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout427_A _07965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13350__A team_01_WB.instance_to_wrap.cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1169_A team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08444__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11397__A2 _07696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09105_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[13\] net664 _05425_
+ _05434_ _05436_ vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_150_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_131_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09036_ _05264_ _05265_ _05302_ _05375_ vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout796_A net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13543__B1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold340 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[126\] vssd1 vssd1 vccd1 vccd1
+ net1875 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold351 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net1886 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1124_X net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold362 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1897 sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1908 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold384 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1919 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold395 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1930 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout963_A _04653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09706__C net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout820 _04632_ vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout831 net834 vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10109__B1 _04678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09938_ _06267_ _06272_ _06277_ vssd1 vssd1 vccd1 vccd1 _06278_ sky130_fd_sc_hd__or3_2
Xfanout842 _03734_ vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__clkbuf_4
Xfanout853 net868 vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__clkbuf_4
Xfanout864 net867 vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__buf_2
Xfanout875 net876 vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09514__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11029__B net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09869_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[12\] net775 _06200_
+ _06201_ _06208_ vssd1 vssd1 vccd1 vccd1 _06209_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout751_X net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout897 _04793_ vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__buf_4
Xhold1040 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2575 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout849_X net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1051 _03452_ vssd1 vssd1 vccd1 vccd1 net2586 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1062 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[57\] vssd1 vssd1 vccd1 vccd1
+ net2597 sky130_fd_sc_hd__dlygate4sd3_1
X_11900_ net2674 net272 net481 vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1073 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 net2608
+ sky130_fd_sc_hd__dlygate4sd3_1
X_12880_ _05779_ net577 net360 vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_29_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1084 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1095 _02093_ vssd1 vssd1 vccd1 vccd1 net2630 sky130_fd_sc_hd__dlygate4sd3_1
X_11831_ net3134 net212 net487 vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__mux2_1
XANTENNA__09278__A1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08338__B net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15740__A net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14550_ net1401 vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__inv_2
X_11762_ net2162 net217 net496 vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__mux2_1
XANTENNA__12821__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ net185 _03959_ _03960_ net723 vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__a211o_1
X_10713_ net557 _07035_ _07052_ vssd1 vssd1 vccd1 vccd1 _07053_ sky130_fd_sc_hd__o21ba_1
XANTENNA__12575__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ net1367 vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11693_ _07889_ _07891_ net614 vssd1 vssd1 vccd1 vccd1 _07892_ sky130_fd_sc_hd__mux2_2
XFILLER_0_82_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16220_ clknet_leaf_139_wb_clk_i net2143 _00208_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__dfrtp_1
X_17951__1466 vssd1 vssd1 vccd1 vccd1 _17951__1466/HI net1466 sky130_fd_sc_hd__conb_1
X_13432_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\]
+ net595 vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__and3_1
XFILLER_0_125_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10644_ _06982_ _06983_ net538 vssd1 vssd1 vccd1 vccd1 _06984_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16151_ clknet_leaf_128_wb_clk_i net2684 _00139_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10575_ _06910_ _06913_ vssd1 vssd1 vccd1 vccd1 _06915_ sky130_fd_sc_hd__or2_2
XANTENNA__10596__A0 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13363_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[11\] _03833_ net827 vssd1 vssd1
+ vccd1 vccd1 _01879_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15102_ net1316 vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__inv_2
X_12314_ net2788 net283 net434 vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16082_ clknet_leaf_131_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[4\]
+ _00070_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13294_ net1069 _07710_ team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1 vccd1
+ vccd1 _03780_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_133_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17642__CLK clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11919__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15033_ net1237 vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__inv_2
X_12245_ net2462 net287 net442 vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__mux2_1
XANTENNA__12888__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12176_ net1857 net253 net448 vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_48 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09753__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08520__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08961__B1 _05266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11127_ _07301_ _07452_ net540 vssd1 vssd1 vccd1 vccd1 _07467_ sky130_fd_sc_hd__mux2_1
X_16984_ clknet_leaf_49_wb_clk_i _02671_ _00967_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11058_ _07381_ _07384_ _07397_ vssd1 vssd1 vccd1 vccd1 _07398_ sky130_fd_sc_hd__and3_1
X_15935_ net1412 vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_60_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10009_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[1\] net775 _06347_ _06348_
+ vssd1 vssd1 vccd1 vccd1 _06349_ sky130_fd_sc_hd__a211o_1
X_15866_ net1202 vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__inv_2
XANTENNA__10520__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08529__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17605_ clknet_leaf_86_wb_clk_i _03292_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_14817_ net1280 vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__inv_2
X_15797_ net1231 vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__inv_2
XFILLER_0_147_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17536_ clknet_leaf_39_wb_clk_i _03223_ _01519_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_14748_ net1187 vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_48_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_80_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12485__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17467_ clknet_leaf_71_wb_clk_i _03154_ _01450_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14679_ net1226 vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__inv_2
XANTENNA__08492__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16418_ clknet_leaf_138_wb_clk_i _02172_ _00401_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17398_ clknet_leaf_12_wb_clk_i _03085_ _01381_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16349_ clknet_leaf_120_wb_clk_i _02103_ _00332_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[72\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09441__A1 _05780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10051__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09992__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18019_ net637 vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11829__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12879__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09095__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09744__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07984_ team_01_WB.instance_to_wrap.cpu.f0.i\[12\] vssd1 vssd1 vccd1 vccd1 _04482_
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_35_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09723_ _06052_ _06054_ _06059_ _06062_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_87_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_87_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09654_ _05983_ _05985_ _05990_ _05993_ vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__or4_4
XANTENNA__10511__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09034__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08605_ net1168 _04846_ _04845_ vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__a21oi_2
X_09585_ _05921_ _05922_ _05923_ _05924_ vssd1 vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout544_A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15560__A net1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11067__B2 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08536_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[18\] net674 _04859_
+ _04867_ _04869_ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12803__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10200__C net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10814__A1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10908__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout332_X net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12395__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08467_ net1001 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[23\] net891
+ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1074_X net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout809_A net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire506 _06463_ vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__clkbuf_2
X_08398_ _04712_ _04737_ _04731_ _04715_ vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_150_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10360_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[17\] net806 net756 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _06700_ sky130_fd_sc_hd__a22o_1
XANTENNA__09557__X _05897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08461__X _04801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09983__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout799_X net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09019_ net1100 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[9\] net893 vssd1
+ vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__and3_1
X_10291_ net990 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[19\] net984 vssd1
+ vssd1 vccd1 vccd1 _06631_ sky130_fd_sc_hd__and3_1
X_12030_ net2319 net211 net463 vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__mux2_1
Xhold170 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[29\] vssd1 vssd1 vccd1 vccd1
+ net1705 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold181 _02028_ vssd1 vssd1 vccd1 vccd1 net1716 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1727 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11542__A2 team_01_WB.instance_to_wrap.cpu.DM0.ihit vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout650 _04821_ vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__buf_6
Xfanout661 _04811_ vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__buf_6
Xfanout672 _04794_ vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__clkbuf_8
Xfanout683 _04783_ vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__buf_8
X_13981_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[0\] _04265_ _04269_ vssd1 vssd1
+ vccd1 vccd1 _04273_ sky130_fd_sc_hd__a21o_1
Xfanout694 net695 vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__clkbuf_8
XANTENNA__17723__Q team_01_WB.instance_to_wrap.cpu.RU0.state\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15720_ net1385 vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__inv_2
XANTENNA__13255__A team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12932_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[13\] net1038 vssd1 vssd1 vccd1
+ vccd1 _03698_ sky130_fd_sc_hd__or2_1
XANTENNA__08349__A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15651_ net1270 vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__inv_2
X_12863_ net2929 net320 net381 vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_122_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09171__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ net1358 vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__inv_2
X_11814_ net2130 net281 net492 vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__mux2_1
X_15582_ net1345 vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__inv_2
X_12794_ net1773 net639 net607 _03624_ vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17321_ clknet_leaf_41_wb_clk_i _03008_ _01304_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10805__A1 _05657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14533_ net1412 vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__inv_2
XANTENNA__10805__B2 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11745_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\]
+ vssd1 vssd1 vccd1 vccd1 _07934_ sky130_fd_sc_hd__xor2_1
XFILLER_0_138_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17252_ clknet_leaf_84_wb_clk_i _02939_ _01235_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_14464_ net1359 vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__inv_2
X_11676_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[16\] _07541_ net715 vssd1 vssd1
+ vccd1 vccd1 _07878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16203_ clknet_leaf_158_wb_clk_i _01963_ _00191_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16074__Q team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13415_ _03874_ _03875_ _03873_ vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_52_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08515__C net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17183_ clknet_leaf_43_wb_clk_i _02870_ _01166_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10627_ net519 net503 vssd1 vssd1 vccd1 vccd1 _06967_ sky130_fd_sc_hd__nand2_2
XFILLER_0_148_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14395_ net1186 vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10033__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16134_ clknet_leaf_157_wb_clk_i _00008_ _00122_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.curr_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__09908__A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13346_ team_01_WB.instance_to_wrap.cpu.f0.i\[11\] net1071 _07677_ team_01_WB.instance_to_wrap.cpu.f0.i\[12\]
+ vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__a31o_1
XANTENNA__09974__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10558_ _04707_ _05151_ net533 vssd1 vssd1 vccd1 vccd1 _06898_ sky130_fd_sc_hd__or3_1
XANTENNA__08371__X _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16065_ clknet_leaf_155_wb_clk_i _01858_ _00053_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\]
+ sky130_fd_sc_hd__dfrtp_4
X_13277_ team_01_WB.instance_to_wrap.cpu.f0.i\[26\] _03747_ vssd1 vssd1 vccd1 vccd1
+ _03766_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10489_ _06826_ _06828_ _05839_ vssd1 vssd1 vccd1 vccd1 _06829_ sky130_fd_sc_hd__a21o_1
X_15016_ net1385 vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__inv_2
X_12228_ net2693 net218 net441 vssd1 vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_121_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11533__A2 net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12159_ net1991 net223 net447 vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17633__Q team_01_WB.instance_to_wrap.cpu.IG0.Instr\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16967_ clknet_leaf_100_wb_clk_i _02654_ _00950_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_15918_ net1415 vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__inv_2
X_16898_ clknet_leaf_56_wb_clk_i _02585_ _00881_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09081__C net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15849_ net1334 vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09789__S net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09370_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[26\] net689 net682 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16562__CLK clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08321_ net992 net954 vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17519_ clknet_leaf_33_wb_clk_i _03206_ _01502_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13994__B1 _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08252_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[29\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[21\]
+ net1051 vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__mux2_1
XANTENNA__10272__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08183_ net2992 net2838 net1052 vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14724__A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10024__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11221__A1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09965__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08722__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1034_A team_01_WB.instance_to_wrap.cpu.RU0.InstrRead vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09717__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_15__f_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09256__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout494_A _07944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13774__S _04146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15555__A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1201_A net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12898__B net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17950__1465 vssd1 vssd1 vccd1 vccd1 _17950__1465/HI net1465 sky130_fd_sc_hd__conb_1
X_07967_ team_01_WB.instance_to_wrap.cpu.f0.i\[31\] vssd1 vssd1 vccd1 vccd1 _04465_
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_71_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout759_A net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09706_ net1154 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[21\] net955
+ vssd1 vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__and3_1
XFILLER_0_156_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_143_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08153__A1 team_01_WB.instance_to_wrap.cpu.f0.read_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09350__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11307__B _05116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09637_ net1136 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[23\] net977
+ vssd1 vssd1 vccd1 vccd1 _05977_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout926_A net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09568_ net1149 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[25\] net971
+ vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13985__B1 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08519_ net1000 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[18\] net935 vssd1
+ vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__and3_1
X_09499_ _05837_ _05838_ vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout714_X net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11323__A team_01_WB.instance_to_wrap.cpu.DM0.data_i\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11530_ net1710 net1171 net588 net1118 vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__a22o_1
XANTENNA__11460__A1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_137_Right_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11042__B _06250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14056__D _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12853__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_122_Left_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11461_ net1169 _04713_ _04753_ vssd1 vssd1 vccd1 vccd1 _07757_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_68_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13201__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13200_ net8 net836 net629 net1701 vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__o22a_1
XFILLER_0_150_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10412_ net1132 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[27\] net977
+ vssd1 vssd1 vccd1 vccd1 _06752_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_78_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10015__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14180_ net1426 _04451_ _04452_ vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__nor3_1
X_11392_ _07697_ _07715_ _04466_ vssd1 vssd1 vccd1 vccd1 _07719_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08632__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13131_ net1607 net851 net632 team_01_WB.instance_to_wrap.a1.ADR_I\[12\] vssd1 vssd1
+ vccd1 vccd1 _02010_ sky130_fd_sc_hd__a22o_1
XANTENNA__16271__D net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12960__A1 _05258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10343_ net1137 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[17\] net946
+ vssd1 vssd1 vccd1 vccd1 _06683_ sky130_fd_sc_hd__and3_1
XFILLER_0_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input55_A wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13062_ net2647 net2637 net852 vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__mux2_1
X_10274_ net1128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[19\] net963
+ vssd1 vssd1 vccd1 vccd1 _06614_ sky130_fd_sc_hd__and3_1
XANTENNA__09166__C net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12013_ net2990 net228 net467 vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__mux2_1
X_17870_ clknet_leaf_129_wb_clk_i _03545_ _01810_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1401 net1402 vssd1 vssd1 vccd1 vccd1 net1401 sky130_fd_sc_hd__buf_4
Xfanout1412 net1414 vssd1 vssd1 vccd1 vccd1 net1412 sky130_fd_sc_hd__buf_4
Xfanout1423 net1424 vssd1 vssd1 vccd1 vccd1 net1423 sky130_fd_sc_hd__buf_4
XFILLER_0_100_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08392__A1 net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16821_ clknet_leaf_118_wb_clk_i _02508_ _00804_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_131_Left_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout480 _07949_ vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__buf_4
Xfanout491 _07944_ vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__buf_8
XANTENNA__11279__A1 _07042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16752_ clknet_leaf_148_wb_clk_i _02439_ _00735_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13964_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[4\]
+ _04220_ _04228_ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__and4_4
XANTENNA__16585__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08144__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15703_ net1216 vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__inv_2
XANTENNA__16069__Q team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12915_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[18\] net1040 vssd1 vssd1 vccd1
+ vccd1 _03686_ sky130_fd_sc_hd__or2_1
X_16683_ clknet_leaf_7_wb_clk_i _02370_ _00666_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08695__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13895_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[0\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[1\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[2\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_17_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11932__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15634_ net1290 vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12846_ net2909 net238 net379 vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__mux2_1
XANTENNA__08366__X _04706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08807__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15565_ net1266 vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__inv_2
XANTENNA__13432__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12777_ net1032 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[17\] vssd1 vssd1 vccd1
+ vccd1 _03613_ sky130_fd_sc_hd__or2_1
X_17304_ clknet_leaf_27_wb_clk_i _02991_ _01287_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14516_ net1407 vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_140_Left_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11451__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11728_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] _07798_ vssd1 vssd1 vccd1
+ vccd1 _07920_ sky130_fd_sc_hd__or2_1
X_15496_ net1375 vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17235_ clknet_leaf_23_wb_clk_i _02922_ _01218_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14447_ net1225 vssd1 vssd1 vccd1 vccd1 _00241_ sky130_fd_sc_hd__inv_2
X_11659_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] _07813_ vssd1 vssd1
+ vccd1 vccd1 _07865_ sky130_fd_sc_hd__or2_1
XANTENNA__18016__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10006__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17166_ clknet_leaf_36_wb_clk_i _02853_ _01149_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09638__A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14378_ net1208 vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__inv_2
XANTENNA__17628__Q team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold906 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2441 sky130_fd_sc_hd__dlygate4sd3_1
X_16117_ clknet_leaf_136_wb_clk_i _01892_ _00105_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[24\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold917 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2452 sky130_fd_sc_hd__dlygate4sd3_1
X_13329_ net564 _07704_ _07733_ net828 vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__a31o_1
XANTENNA__12951__B2 _03710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold928 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold939 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2474 sky130_fd_sc_hd__dlygate4sd3_1
X_17097_ clknet_leaf_39_wb_clk_i _02784_ _01080_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14153__B1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16048_ clknet_leaf_148_wb_clk_i _01841_ _00036_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_122_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11506__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08870_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[3\] net649 _05193_ _05197_
+ _05207_ vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_32_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1606 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net3141 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09580__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1617 net107 vssd1 vssd1 vccd1 vccd1 net3152 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1628 team_01_WB.instance_to_wrap.cpu.DM0.state\[2\] vssd1 vssd1 vccd1 vccd1 net3163
+ sky130_fd_sc_hd__dlygate4sd3_1
X_17999_ net635 vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__clkbuf_1
Xhold1639 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 net3174
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12003__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11842__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13182__X _03738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09422_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[28\] net686 net669 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__a22o_1
XANTENNA__11690__A1 _07553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08717__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09353_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[25\] net673 net659 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[25\]
+ _05683_ vssd1 vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__a221o_1
XANTENNA__08436__B net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08304_ net990 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[30\] net972 vssd1
+ vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__and3_1
XANTENNA__10245__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09284_ net1009 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[22\] net896 vssd1
+ vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08235_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[46\] net2585 net1042 vssd1 vssd1
+ vccd1 vccd1 _03452_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12673__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1151_A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout507_A _06098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09399__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08166_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[115\] net1748 net1054 vssd1 vssd1
+ vccd1 vccd1 _03521_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12942__A1 _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08097_ _04564_ _04565_ _04566_ _04567_ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__or4_1
XFILLER_0_31_857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08610__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1416_A net1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1037_X net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload90 clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload90/Y sky130_fd_sc_hd__inv_6
XANTENNA__14144__B1 _04245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13498__A2 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout497_X net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout876_A net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09283__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout664_X net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08999_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] net595 vssd1 vssd1 vccd1
+ vccd1 _05339_ sky130_fd_sc_hd__nand2_1
XANTENNA__09323__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_117_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_117_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout831_X net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10961_ net546 _06438_ _06939_ vssd1 vssd1 vccd1 vccd1 _07301_ sky130_fd_sc_hd__o21ba_1
XANTENNA__12848__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13670__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11752__S net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout929_X net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12700_ net1913 net240 net383 vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__mux2_1
X_13680_ team_01_WB.instance_to_wrap.cpu.c0.count\[6\] _04102_ vssd1 vssd1 vccd1 vccd1
+ _04103_ sky130_fd_sc_hd__and2_1
XANTENNA__11681__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10892_ net562 _07208_ _07209_ _07230_ vssd1 vssd1 vccd1 vccd1 _07232_ sky130_fd_sc_hd__a31o_1
XFILLER_0_35_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12631_ net2249 net202 net394 vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08346__B net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10236__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15350_ net1256 vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12562_ net2638 net206 net401 vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14301_ net1328 vssd1 vssd1 vccd1 vccd1 _00095_ sky130_fd_sc_hd__inv_2
X_11513_ net1558 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[5\] net877 vssd1 vssd1
+ vccd1 vccd1 _03336_ sky130_fd_sc_hd__mux2_1
X_15281_ net1397 vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__inv_2
XANTENNA__12583__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14364__A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12493_ net2926 net215 net409 vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_117_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17020_ clknet_leaf_50_wb_clk_i _02707_ _01003_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_117_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14232_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[0\] vssd1 vssd1 vccd1
+ vccd1 _02255_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_22_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09929__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11444_ _07675_ net325 _07746_ vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__and3b_1
XFILLER_0_34_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12933__A1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14163_ net1426 _04442_ vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__nor2_1
X_11375_ _07703_ vssd1 vssd1 vccd1 vccd1 _07704_ sky130_fd_sc_hd__inv_2
XANTENNA__10944__A0 _06495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08601__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13114_ net96 net844 net634 net1598 vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__a22o_1
XANTENNA__14135__B1 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10326_ net1129 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[18\] net972
+ vssd1 vssd1 vccd1 vccd1 _06666_ sky130_fd_sc_hd__and3_1
X_14094_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[77\] _04235_ _04266_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__a22o_1
XANTENNA__11927__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13045_ net2553 net2444 net865 vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__mux2_1
X_17922_ net1529 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
X_10257_ _06533_ _06568_ _06596_ vssd1 vssd1 vccd1 vccd1 _06597_ sky130_fd_sc_hd__or3_1
XFILLER_0_147_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1220 net1221 vssd1 vssd1 vccd1 vccd1 net1220 sky130_fd_sc_hd__buf_4
Xfanout1231 net1232 vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__buf_4
XANTENNA__13427__B _04971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10188_ _04750_ _05006_ _05376_ vssd1 vssd1 vccd1 vccd1 _06528_ sky130_fd_sc_hd__nand3_1
Xfanout1242 net1304 vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__buf_2
X_17853_ clknet_leaf_96_wb_clk_i net1783 _01793_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[123\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1253 net1255 vssd1 vssd1 vccd1 vccd1 net1253 sky130_fd_sc_hd__buf_4
Xfanout1264 net1269 vssd1 vssd1 vccd1 vccd1 net1264 sky130_fd_sc_hd__buf_2
X_16804_ clknet_leaf_84_wb_clk_i _02491_ _00787_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1275 net1277 vssd1 vssd1 vccd1 vccd1 net1275 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_4_14__f_wb_clk_i_X clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1286 net1289 vssd1 vssd1 vccd1 vccd1 net1286 sky130_fd_sc_hd__buf_4
Xfanout1297 net1298 vssd1 vssd1 vccd1 vccd1 net1297 sky130_fd_sc_hd__buf_4
X_17784_ clknet_leaf_117_wb_clk_i net2738 _01724_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14996_ net1379 vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__inv_2
X_16735_ clknet_leaf_42_wb_clk_i _02422_ _00718_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13947_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[3\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__and2_2
XANTENNA__12758__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14539__A net1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11662__S net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16666_ clknet_leaf_78_wb_clk_i _02353_ _00649_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11672__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13878_ team_01_WB.instance_to_wrap.cpu.RU0.state\[0\] _03579_ _04136_ vssd1 vssd1
+ vccd1 vccd1 _00006_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15617_ net1282 vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__inv_2
X_12829_ net1035 _07476_ net365 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\]
+ net1063 vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__a32o_1
X_16597_ clknet_leaf_114_wb_clk_i _02284_ _00580_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13413__A2 _05116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15548_ net1252 vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15479_ net1244 vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__inv_2
XANTENNA__12493__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08840__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08020_ team_01_WB.instance_to_wrap.cpu.K0.keyvalid _04515_ vssd1 vssd1 vccd1 vccd1
+ _04516_ sky130_fd_sc_hd__nand2_2
XFILLER_0_141_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17218_ clknet_leaf_57_wb_clk_i _02905_ _01201_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold703 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[17\] vssd1 vssd1 vccd1 vccd1
+ net2238 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12924__A1 _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11727__A2 _07323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17149_ clknet_leaf_65_wb_clk_i _02836_ _01132_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold714 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2249 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10307__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold725 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2260 sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2271 sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2282 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14126__B1 _04241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold758 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2293 sky130_fd_sc_hd__dlygate4sd3_1
X_09971_ _06303_ _06304_ _06309_ _06310_ vssd1 vssd1 vccd1 vccd1 _06311_ sky130_fd_sc_hd__or4_2
Xhold769 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[18\] vssd1 vssd1 vccd1 vccd1
+ net2304 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11837__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08922_ net531 net521 vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_90_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08853_ net1109 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[3\] net884 vssd1
+ vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__and3_1
Xhold1403 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2938 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09534__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout192_A _07634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1414 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[70\] vssd1 vssd1 vccd1 vccd1
+ net2949 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1425 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[118\] vssd1 vssd1 vccd1 vccd1
+ net2960 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1436 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2971 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1447 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2982 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10042__A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08784_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[0\] net664 _05121_ _05122_
+ _05123_ vssd1 vssd1 vccd1 vccd1 _05124_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13637__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1458 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2993 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_140_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1469 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net3004 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12668__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08659__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13652__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout457_A _07956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1199_A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10466__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09320__A3 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09405_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[27\] net686 net684 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout624_A _04628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10218__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09336_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[24\] net689 net682 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[24\]
+ _05662_ vssd1 vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__a221o_1
XANTENNA__08734__X _05074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout412_X net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09267_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[20\] net696 net660 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[20\]
+ _05606_ vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1154_X net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11601__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08218_ net2894 net2828 net1047 vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__mux2_1
X_09198_ net1087 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[17\] net888
+ vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout993_A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08149_ _04610_ _04611_ _04615_ _04618_ vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_43_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1321_X net1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14912__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11160_ net334 net337 _07383_ vssd1 vssd1 vccd1 vccd1 _07500_ sky130_fd_sc_hd__mux2_1
XANTENNA__10500__A_N net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout781_X net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11747__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout879_X net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10111_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[6\] _04649_ net738 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06451_ sky130_fd_sc_hd__a22o_1
X_11091_ _06858_ _06882_ _07412_ _07430_ vssd1 vssd1 vccd1 vccd1 _07431_ sky130_fd_sc_hd__o211a_1
X_10042_ net994 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[0\] net958 vssd1
+ vssd1 vccd1 vccd1 _06382_ sky130_fd_sc_hd__and3_1
XANTENNA__09544__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold30 team_01_WB.instance_to_wrap.cpu.f0.write_data\[10\] vssd1 vssd1 vccd1 vccd1
+ net1565 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09444__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold41 _02011_ vssd1 vssd1 vccd1 vccd1 net1576 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[23\] vssd1 vssd1 vccd1 vccd1 net1587
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14850_ net1346 vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__inv_2
Xhold63 team_01_WB.instance_to_wrap.a1.ADR_I\[29\] vssd1 vssd1 vccd1 vccd1 net1598
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[26\] vssd1 vssd1 vccd1 vccd1 net1609
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 team_01_WB.instance_to_wrap.a1.ADR_I\[0\] vssd1 vssd1 vccd1 vccd1 net1620
+ sky130_fd_sc_hd__dlygate4sd3_1
X_13801_ _01835_ _04173_ vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__nand2_1
Xhold96 _02008_ vssd1 vssd1 vccd1 vccd1 net1631 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09741__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12578__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input18_A DAT_I[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14781_ net1236 vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__inv_2
XANTENNA__09847__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[13\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17731__Q team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11993_ net2499 net191 net467 vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__mux2_1
X_16520_ clknet_leaf_1_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[18\]
+ _00503_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13732_ _04507_ team_01_WB.instance_to_wrap.a1.READ_I team_01_WB.instance_to_wrap.a1.curr_state\[0\]
+ _04509_ team_01_WB.instance_to_wrap.a1.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 _00009_
+ sky130_fd_sc_hd__a32o_1
X_10944_ _06495_ _06526_ net339 _06562_ net550 net539 vssd1 vssd1 vccd1 vccd1 _07284_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10457__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16451_ clknet_leaf_72_wb_clk_i _02205_ _00434_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13663_ _07639_ _04093_ _04094_ net728 vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__a211o_1
XFILLER_0_128_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10875_ _07024_ _07214_ net514 vssd1 vssd1 vccd1 vccd1 _07215_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15402_ net1284 vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__inv_2
X_12614_ net3110 net297 net398 vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10209__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11406__A1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16382_ clknet_leaf_88_wb_clk_i _02136_ _00365_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[105\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09075__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11214__C _07251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13594_ net198 net194 _07810_ _07887_ net644 vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__o2111a_1
Xclkbuf_leaf_85_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15333_ net1263 vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__inv_2
X_12545_ net2732 net282 net405 vssd1 vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_54_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15264_ net1278 vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__inv_2
X_12476_ net2650 net285 net414 vssd1 vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__mux2_1
X_17003_ clknet_leaf_8_wb_clk_i _02690_ _00986_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_14215_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[17\] vssd1 vssd1 vccd1
+ vccd1 _02272_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08523__C net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_5 _03654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11427_ _04480_ _07738_ _07699_ _07689_ vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__a211oi_1
X_15195_ net1255 vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__inv_2
X_14146_ _04424_ _04426_ _04428_ _04430_ vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__or4_1
XANTENNA__09783__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11358_ net1071 _07679_ vssd1 vssd1 vccd1 vccd1 _07687_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10309_ net1130 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[18\] net980
+ vssd1 vssd1 vccd1 vccd1 _06649_ sky130_fd_sc_hd__and3_1
X_14077_ _04358_ _04360_ _04362_ _04364_ vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__or4_1
X_11289_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] _07628_ vssd1 vssd1 vccd1
+ vccd1 _07629_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13028_ net2594 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[66\] net863 vssd1 vssd1
+ vccd1 vccd1 _02097_ sky130_fd_sc_hd__mux2_1
X_17905_ net1440 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
Xfanout1050 net1051 vssd1 vssd1 vccd1 vccd1 net1050 sky130_fd_sc_hd__clkbuf_4
Xfanout1061 team_01_WB.instance_to_wrap.cpu.RU0.state\[5\] vssd1 vssd1 vccd1 vccd1
+ net1061 sky130_fd_sc_hd__buf_4
X_17836_ clknet_leaf_102_wb_clk_i net2944 _01776_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[106\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1072 team_01_WB.instance_to_wrap.cpu.f0.i\[7\] vssd1 vssd1 vccd1 vccd1 net1072
+ sky130_fd_sc_hd__clkbuf_2
Xfanout1083 net1089 vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__buf_2
Xfanout1094 net1096 vssd1 vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__buf_2
XANTENNA__12488__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17641__Q team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17767_ clknet_leaf_98_wb_clk_i _03443_ _01707_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[37\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__12889__B1_N net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13634__A2 _07290_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14979_ net1250 vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16718_ clknet_leaf_36_wb_clk_i _02405_ _00701_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17698_ clknet_leaf_134_wb_clk_i _03382_ _01639_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16649_ clknet_leaf_40_wb_clk_i _02336_ _00632_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09066__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09121_ net1110 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[14\] net941
+ vssd1 vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__and3_1
XANTENNA__08274__A0 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10081__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire961_A _04656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09052_ net1109 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[12\] net890
+ vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08003_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1 vccd1 vccd1
+ _04501_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_133_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold500 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2035 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10037__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold511 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[34\] vssd1 vssd1 vccd1 vccd1
+ net2046 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold522 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2057 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout205_A _07855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold533 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2068 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09826__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13570__A1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09774__B1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold544 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2079 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold555 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2090 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold566 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[1\] vssd1 vssd1 vccd1 vccd1 net2101
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2112 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold588 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2123 sky130_fd_sc_hd__dlygate4sd3_1
X_09954_ net998 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[3\] net957 vssd1
+ vssd1 vccd1 vccd1 _06294_ sky130_fd_sc_hd__and3_1
Xhold599 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2134 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1114_A net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09526__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08905_ net1107 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[2\] net884 vssd1
+ vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__and3_1
X_09885_ net998 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[5\] net974 vssd1
+ vssd1 vccd1 vccd1 _06225_ sky130_fd_sc_hd__and3_1
Xhold1200 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2735 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1211 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[86\] vssd1 vssd1 vccd1 vccd1
+ net2746 sky130_fd_sc_hd__dlygate4sd3_1
X_08836_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[1\] net686 _05158_ _05162_
+ _05171_ vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__a2111o_1
Xhold1222 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[55\] vssd1 vssd1 vccd1 vccd1
+ net2757 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1233 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2768 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1244 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[66\] vssd1 vssd1 vccd1 vccd1
+ net2779 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10203__C _04662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1255 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[63\] vssd1 vssd1 vccd1 vccd1
+ net2790 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09561__A _05898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1266 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[72\] vssd1 vssd1 vccd1 vccd1
+ net2801 sky130_fd_sc_hd__dlygate4sd3_1
X_08767_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[4\] net650 _05082_ _05089_
+ _05090_ vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12398__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1277 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2812 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout362_X net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1288 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2823 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1299 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2834 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout839_A _03734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10439__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08698_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[7\] net690 _05015_ _05023_
+ _05027_ vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_105_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14907__A net1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout627_X net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1369_X net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10660_ _06998_ _06999_ net541 vssd1 vssd1 vccd1 vccd1 _07000_ sky130_fd_sc_hd__mux2_1
XANTENNA__08464__X _04804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14050__A2 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09319_ _04844_ _05570_ _05620_ _05658_ vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_81_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08804__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10591_ net375 _06897_ _06899_ _06904_ vssd1 vssd1 vccd1 vccd1 _06931_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_153_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12330_ net2814 net248 net429 vssd1 vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_153_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout996_X net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08343__C net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12261_ net2606 net219 net437 vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__mux2_1
XANTENNA__12861__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14000_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[1\] _04249_ _04259_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13561__A1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11212_ _07550_ _07551_ _07547_ vssd1 vssd1 vccd1 vccd1 _07552_ sky130_fd_sc_hd__or3b_1
XANTENNA__09736__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12192_ net2268 net222 net443 vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10914__A3 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13258__A team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11143_ _07180_ _07317_ net516 vssd1 vssd1 vccd1 vccd1 _07483_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 ADR_O[0] sky130_fd_sc_hd__buf_2
XANTENNA__13313__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_132_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_132_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 ADR_O[1] sky130_fd_sc_hd__buf_2
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__buf_2
X_11074_ net371 _07223_ _05529_ vssd1 vssd1 vccd1 vccd1 _07414_ sky130_fd_sc_hd__or3b_1
X_15951_ net1412 vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__inv_2
X_14902_ net1247 vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__inv_2
X_10025_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[1\] net766 _06358_ _06364_
+ vssd1 vssd1 vccd1 vccd1 _06365_ sky130_fd_sc_hd__o22a_1
X_15882_ net1347 vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_129_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09471__A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17621_ clknet_leaf_6_wb_clk_i _03306_ _01562_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_14833_ net1423 vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11627__A1 _07588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14764_ net1261 vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__inv_2
X_17552_ clknet_leaf_146_wb_clk_i _03239_ _01535_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12101__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08087__A team_01_WB.instance_to_wrap.cpu.f0.i\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11976_ net2361 net230 net473 vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_38_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13715_ net3104 _04102_ vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__nor2_1
X_16503_ clknet_leaf_2_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[1\]
+ _00486_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08518__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10927_ _06980_ _07227_ _07265_ _06921_ _07185_ vssd1 vssd1 vccd1 vccd1 _07267_ sky130_fd_sc_hd__o221a_1
X_17483_ clknet_leaf_5_wb_clk_i _03170_ _01466_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_14695_ net1210 vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__inv_2
XANTENNA__11940__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16434_ clknet_leaf_133_wb_clk_i _02188_ _00417_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13646_ _03868_ _03880_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10858_ _06158_ net373 _06216_ net340 net550 net539 vssd1 vssd1 vccd1 vccd1 _07198_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_67_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14041__A2 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12938__A2_N _03701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16365_ clknet_leaf_122_wb_clk_i _02119_ _00348_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[88\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13577_ net986 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] _04022_ _04023_
+ vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10789_ _04919_ _07125_ _07128_ vssd1 vssd1 vccd1 vccd1 _07129_ sky130_fd_sc_hd__a21o_1
X_15316_ net1378 vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__inv_2
X_12528_ net2501 net245 net404 vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16296_ clknet_leaf_97_wb_clk_i _02050_ _00279_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15247_ net1386 vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__inv_2
X_12459_ net2502 net220 net413 vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15178_ net1385 vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__inv_2
XANTENNA__09220__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10366__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[17\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08550__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16540__Q team_01_WB.instance_to_wrap.cpu.DM0.data_i\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14129_ _04404_ _04411_ _04413_ _04414_ vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__or4_1
Xfanout309 net310 vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09084__C net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_77_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09670_ net1136 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[22\] net965
+ vssd1 vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__and3_1
X_08621_ _04955_ _04957_ _04958_ _04960_ vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__or4_1
X_17819_ clknet_leaf_93_wb_clk_i net2800 _01759_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[89\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12011__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11618__A1 _07088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08552_ net999 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[19\] net897 vssd1
+ vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__and3_1
XANTENNA__10320__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08483_ net1107 net889 vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__and2_2
XANTENNA__11850__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11703__X _07900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10841__A2 _06636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14032__A2 _04246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1064_A net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09104_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[13\] net695 _05423_
+ _05424_ _05429_ vssd1 vssd1 vccd1 vccd1 _05444_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11151__A _07449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09995__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16032__RESET_B net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09035_ _05338_ _05374_ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__nand2_1
XFILLER_0_142_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12681__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1329_A net1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13543__A1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold330 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1865 sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 _02157_ vssd1 vssd1 vccd1 vccd1 net1876 sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net1887 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout691_A _04772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout789_A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold363 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1898 sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1909 sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1920 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1931 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14099__A2 _04245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout810 _04639_ vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout821 net824 vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__buf_6
X_09937_ _06273_ _06274_ _06276_ vssd1 vssd1 vccd1 vccd1 _06277_ sky130_fd_sc_hd__or3_1
Xfanout832 net834 vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__clkbuf_2
Xfanout843 net851 vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout577_X net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout956_A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout854 net855 vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10419__A_N net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout865 net866 vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13806__A team_01_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout876 net877 vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__buf_2
X_09868_ _06202_ _06203_ _06204_ _06207_ vssd1 vssd1 vccd1 vccd1 _06208_ sky130_fd_sc_hd__or4_1
Xfanout887 _04799_ vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__buf_4
Xfanout898 net899 vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__buf_4
XANTENNA__08459__X _04799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1030 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[75\] vssd1 vssd1 vccd1 vccd1
+ net2565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1041 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2576 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08819_ net1105 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[1\] net907 vssd1
+ vssd1 vccd1 vccd1 _05159_ sky130_fd_sc_hd__and3_1
Xhold1052 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[27\] vssd1 vssd1 vccd1 vccd1
+ net2587 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1063 _02096_ vssd1 vssd1 vccd1 vccd1 net2598 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout744_X net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09799_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[14\] net750 net743 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06139_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_29_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1074 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[96\] vssd1 vssd1 vccd1 vccd1
+ net2609 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1085 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[14\] vssd1 vssd1 vccd1 vccd1
+ net2620 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11609__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1096 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2631 sky130_fd_sc_hd__dlygate4sd3_1
X_11830_ net2558 net214 net489 vssd1 vssd1 vccd1 vccd1 _03147_ sky130_fd_sc_hd__mux2_1
XANTENNA__10230__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12806__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09278__A2 _05615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout911_X net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11085__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11761_ net2248 _07831_ net496 vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__mux2_1
XANTENNA__12856__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11760__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13500_ net196 net192 _07826_ net642 vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_155_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ _06934_ _07043_ _07051_ _06963_ _07048_ vssd1 vssd1 vccd1 vccd1 _07052_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_155_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ net1347 vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__inv_2
X_11692_ _07808_ _07890_ vssd1 vssd1 vccd1 vccd1 _07891_ sky130_fd_sc_hd__nor2_1
XANTENNA__08635__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14023__A2 _04221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13431_ _03890_ _03891_ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10643_ _06671_ _06707_ net544 vssd1 vssd1 vccd1 vccd1 _06983_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10045__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09986__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16150_ clknet_leaf_128_wb_clk_i _01913_ _00138_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11242__C1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13362_ net586 _07684_ _03832_ _03831_ net565 vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__a32o_1
XFILLER_0_51_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10574_ _06910_ _06913_ vssd1 vssd1 vccd1 vccd1 _06914_ sky130_fd_sc_hd__nor2_1
XANTENNA__10596__A1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09450__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15101_ net1240 vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__inv_2
X_12313_ net2004 net249 net434 vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16081_ clknet_leaf_130_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[3\]
+ _00069_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[3\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12591__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13293_ _03746_ _03778_ _04518_ vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_146_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13534__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15032_ net1209 vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__inv_2
X_12244_ net2908 net255 net440 vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__mux2_1
XANTENNA__08370__A team_01_WB.instance_to_wrap.cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11545__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_111_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08801__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12175_ net2980 net257 net449 vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__mux2_1
XANTENNA__10899__A2 _07238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08961__A1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11126_ net535 _06952_ _06954_ _07465_ _05262_ vssd1 vssd1 vccd1 vccd1 _07466_ sky130_fd_sc_hd__o311a_1
XANTENNA__10899__X _07239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16983_ clknet_leaf_16_wb_clk_i _02670_ _00966_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11935__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15934_ net1415 vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__inv_2
X_11057_ _07395_ _07396_ vssd1 vssd1 vccd1 vccd1 _07397_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09910__B1 _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10008_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[1\] net822 net773 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06348_ sky130_fd_sc_hd__a22o_1
X_15865_ net1346 vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__inv_2
XANTENNA__09632__C net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17604_ clknet_leaf_86_wb_clk_i _03291_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_14816_ net1235 vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__inv_2
X_15796_ net1230 vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__inv_2
XANTENNA__09269__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17535_ clknet_leaf_43_wb_clk_i _03222_ _01518_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14747_ net1194 vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__inv_2
X_11959_ net576 _07945_ _07951_ vssd1 vssd1 vccd1 vccd1 _07952_ sky130_fd_sc_hd__and3_4
XANTENNA__14547__A net1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13865__A_N net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18019__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11670__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10284__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17466_ clknet_leaf_78_wb_clk_i _03153_ _01449_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_14678_ net1204 vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_15_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13629_ net989 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] _04066_ _04067_
+ vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__a22o_1
X_16417_ clknet_leaf_126_wb_clk_i _02171_ _00400_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16535__Q team_01_WB.instance_to_wrap.cpu.DM0.data_i\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_17_Left_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17397_ clknet_leaf_110_wb_clk_i _03084_ _01380_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_150_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09977__B1 _04659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16348_ clknet_leaf_97_wb_clk_i _02102_ _00331_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[71\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16279_ clknet_leaf_125_wb_clk_i _02033_ _00262_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_89_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13525__A1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18018_ net1512 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__buf_2
XANTENNA_wire378_X net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08711__C net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16270__Q team_01_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10315__A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12006__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07983_ team_01_WB.instance_to_wrap.cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1 _04481_
+ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_26_Left_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11845__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09722_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[21\] net809 net770 _06060_
+ _06061_ vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11839__A1 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09901__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09653_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[23\] net752 _05991_
+ _05992_ net768 vssd1 vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09542__C net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_157_wb_clk_i_X clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08604_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[15\] net703 _04931_ _04943_
+ vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__o22ai_4
X_09584_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[25\] net809 _05903_
+ _05906_ _05909_ vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_54_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08535_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[18\] net664 _04852_
+ _04858_ _04866_ vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12676__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08466_ net1006 net892 vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__and2_4
XPHY_EDGE_ROW_35_Left_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08455__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14005__A2 _04221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09680__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13213__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout704_A _04758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08397_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] net712 net709 vssd1 vssd1
+ vccd1 vccd1 _04737_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1067_X net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09968__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09432__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09018_ net1100 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[9\] net898 vssd1
+ vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__and3_1
XANTENNA__09286__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13516__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10290_ net1134 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[19\] net968
+ vssd1 vssd1 vccd1 vccd1 _06630_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout694_X net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12724__C1 net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold160 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1695 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 net121 vssd1 vssd1 vccd1 vccd1 net1706 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10225__A _05338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold182 net93 vssd1 vssd1 vccd1 vccd1 net1717 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[2\] vssd1 vssd1 vccd1 vccd1
+ net1728 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout640 _03572_ vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout959_X net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout651 _04821_ vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13095__X _03719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11755__S net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout662 _04808_ vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__clkbuf_8
X_13980_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[48\] _04236_ _04259_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__a22o_1
Xfanout673 _04794_ vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__clkbuf_4
Xfanout684 _04780_ vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__clkbuf_8
Xfanout695 _04768_ vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_126_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12931_ net584 _07757_ _03694_ vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12862_ net2865 net307 net381 vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__mux2_1
X_15650_ net1319 vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_122_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ net2604 net252 net494 vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__mux2_1
X_14601_ net1358 vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__inv_2
X_15581_ net1236 vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__inv_2
XANTENNA__12586__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10895__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12793_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] net1061 net362 _03623_
+ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14532_ net1421 vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__inv_2
X_17320_ clknet_leaf_63_wb_clk_i _03007_ _01303_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10805__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11744_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[3\] net716 net615 vssd1 vssd1
+ vccd1 vccd1 _07933_ sky130_fd_sc_hd__o21a_1
XFILLER_0_28_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14463_ net1225 vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__inv_2
XANTENNA__11503__B _07756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17251_ clknet_leaf_63_wb_clk_i _02938_ _01234_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11675_ net2559 net267 net502 vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__mux2_1
XANTENNA__09959__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16202_ clknet_leaf_159_wb_clk_i _01962_ _00190_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13414_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] _05224_ vssd1 vssd1 vccd1
+ vccd1 _03875_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17182_ clknet_leaf_80_wb_clk_i _02869_ _01165_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10626_ net553 _06965_ vssd1 vssd1 vccd1 vccd1 _06966_ sky130_fd_sc_hd__and2_1
X_14394_ net1189 vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09423__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16133_ clknet_leaf_126_wb_clk_i _00024_ _00121_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.state\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_153_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13345_ _04482_ _07678_ vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__nand2_1
X_10557_ net545 net533 _06858_ vssd1 vssd1 vccd1 vccd1 _06897_ sky130_fd_sc_hd__or3_1
XANTENNA__13507__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16064_ clknet_leaf_155_wb_clk_i _01857_ _00052_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\]
+ sky130_fd_sc_hd__dfrtp_4
X_13276_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[29\] net825 _07650_ _03765_
+ vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__o22a_1
X_10488_ _06750_ _06819_ _06823_ _06827_ _05902_ vssd1 vssd1 vccd1 vccd1 _06828_ sky130_fd_sc_hd__a2111o_1
X_15015_ net1396 vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12227_ net2013 net222 net439 vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__mux2_1
XANTENNA__09924__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12158_ net2469 net191 net447 vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__mux2_1
XANTENNA__11665__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11109_ net344 _06409_ _07439_ _07448_ vssd1 vssd1 vccd1 vccd1 _07449_ sky130_fd_sc_hd__o31a_2
X_16966_ clknet_leaf_91_wb_clk_i _02653_ _00949_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12089_ net2951 net314 net461 vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15917_ net1417 vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__inv_2
X_16897_ clknet_leaf_54_wb_clk_i _02584_ _00880_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15848_ net1334 vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12496__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15779_ net1206 vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_914 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08320_ net1159 net1166 net1165 net1162 vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__and4bb_4
XFILLER_0_115_86 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17518_ clknet_leaf_28_wb_clk_i _03205_ _01501_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08706__C net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08251_ net2797 net3033 net1042 vssd1 vssd1 vccd1 vccd1 _03436_ sky130_fd_sc_hd__mux2_1
X_17449_ clknet_leaf_36_wb_clk_i _03136_ _01432_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08182_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[99\] net2236 net1054 vssd1 vssd1
+ vccd1 vccd1 _03505_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09414__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08622__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09537__C net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08441__C net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10980__B2 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12812__X _03637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout487_A _07947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09705_ net997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[21\] net952 vssd1
+ vssd1 vccd1 vccd1 _06045_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout654_A _04817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1396_A net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09636_ net1135 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[23\] net981
+ vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_43_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09567_ net997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[25\] net970 vssd1
+ vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout821_A net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout442_X net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout919_A net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12788__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08518_ net1001 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[18\] net883 vssd1
+ vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__and3_1
X_09498_ _04706_ _05836_ vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__or2_1
XANTENNA__09653__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08449_ net1112 net902 vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__and2_1
XANTENNA__11323__B team_01_WB.instance_to_wrap.cpu.DM0.data_i\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout707_X net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14915__A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11460_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] _04713_ net718 _04751_ vssd1
+ vssd1 vccd1 vccd1 _07756_ sky130_fd_sc_hd__o22a_4
XFILLER_0_92_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09405__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10411_ net1131 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[27\] net958
+ vssd1 vssd1 vccd1 vccd1 _06751_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11391_ team_01_WB.instance_to_wrap.cpu.f0.i\[30\] _07716_ _07717_ vssd1 vssd1 vccd1
+ vccd1 _03393_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_78_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08613__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13130_ net1575 net843 net631 team_01_WB.instance_to_wrap.a1.ADR_I\[13\] vssd1 vssd1
+ vccd1 vccd1 _02011_ sky130_fd_sc_hd__a22o_1
X_10342_ net1137 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[17\] net968
+ vssd1 vssd1 vccd1 vccd1 _06682_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10971__A1 _06920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10971__B2 _06928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13061_ net2205 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[33\] net865 vssd1 vssd1
+ vccd1 vccd1 _02064_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10273_ net1128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[19\] net958
+ vssd1 vssd1 vccd1 vccd1 _06613_ sky130_fd_sc_hd__and3_1
XFILLER_0_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12012_ net2972 net286 net469 vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__mux2_1
XANTENNA_input48_A wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1402 net1409 vssd1 vssd1 vccd1 vccd1 net1402 sky130_fd_sc_hd__buf_4
Xfanout1413 net1414 vssd1 vssd1 vccd1 vccd1 net1413 sky130_fd_sc_hd__buf_4
XANTENNA__17734__Q team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout1424 net1425 vssd1 vssd1 vccd1 vccd1 net1424 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_39_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16820_ clknet_leaf_66_wb_clk_i _02507_ _00803_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_6_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout470 _07953_ vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__buf_8
Xfanout481 _07949_ vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__buf_6
Xfanout492 _07944_ vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__buf_4
X_16751_ clknet_leaf_34_wb_clk_i _02438_ _00734_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13963_ _04231_ _04237_ _04239_ vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__and3_4
XANTENNA__09341__A1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15702_ net1256 vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__inv_2
X_12914_ net360 _03684_ net1036 vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__o21ai_1
X_13894_ _04140_ net572 _04198_ vssd1 vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__and3_1
X_16682_ clknet_leaf_9_wb_clk_i _02369_ _00665_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_15633_ net1420 vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__inv_2
X_12845_ net2283 net269 net379 vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10239__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15564_ net1259 vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12776_ net1032 _07231_ vssd1 vssd1 vccd1 vccd1 _03612_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09644__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17303_ clknet_leaf_16_wb_clk_i _02990_ _01286_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08526__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14515_ net1415 vssd1 vssd1 vccd1 vccd1 _00309_ sky130_fd_sc_hd__inv_2
XANTENNA__11233__B _07265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11727_ net718 _07323_ net615 _07918_ vssd1 vssd1 vccd1 vccd1 _07919_ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_3_0_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15495_ net1390 vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17234_ clknet_leaf_110_wb_clk_i _02921_ _01217_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11658_ net719 _07171_ net616 _07863_ vssd1 vssd1 vccd1 vccd1 _07864_ sky130_fd_sc_hd__o211a_1
X_14446_ net1307 vssd1 vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10609_ _06438_ net372 net546 vssd1 vssd1 vccd1 vccd1 _06949_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12400__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14377_ net1208 vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__inv_2
X_17165_ clknet_leaf_107_wb_clk_i _02852_ _01148_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11589_ _07805_ vssd1 vssd1 vccd1 vccd1 _07806_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold907 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2442 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13328_ team_01_WB.instance_to_wrap.cpu.f0.i\[16\] _03743_ _03801_ net587 vssd1 vssd1
+ vccd1 vccd1 _03806_ sky130_fd_sc_hd__o211a_1
X_16116_ clknet_leaf_136_wb_clk_i _01891_ _00104_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[23\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold918 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2453 sky130_fd_sc_hd__dlygate4sd3_1
Xhold929 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2464 sky130_fd_sc_hd__dlygate4sd3_1
X_17096_ clknet_leaf_61_wb_clk_i _02783_ _01079_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13259_ team_01_WB.instance_to_wrap.cpu.f0.i\[23\] net1069 _07710_ vssd1 vssd1 vccd1
+ vccd1 _03751_ sky130_fd_sc_hd__or3_1
XFILLER_0_0_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16047_ clknet_leaf_150_wb_clk_i _01840_ _00035_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__17644__Q team_01_WB.instance_to_wrap.cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1607 team_01_WB.instance_to_wrap.cpu.K0.code\[3\] vssd1 vssd1 vccd1 vccd1 net3142
+ sky130_fd_sc_hd__dlygate4sd3_1
X_17998_ net636 vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__clkbuf_1
Xhold1618 team_01_WB.instance_to_wrap.a1.curr_state\[0\] vssd1 vssd1 vccd1 vccd1 net3153
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1629 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net3164 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09092__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16949_ clknet_leaf_118_wb_clk_i _02636_ _00932_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10031__C net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09421_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[28\] net657 net652 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09352_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[25\] net660 net657 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[25\]
+ _05684_ vssd1 vssd1 vccd1 vccd1 _05692_ sky130_fd_sc_hd__a221o_1
X_08303_ net992 net972 vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__and2_4
X_09283_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[22\] net922
+ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__and3_1
XANTENNA__12954__S net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout235_A net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10650__A0 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08234_ net2774 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[39\] net1048 vssd1 vssd1
+ vccd1 vccd1 _03453_ sky130_fd_sc_hd__mux2_1
XANTENNA__08292__X _04632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13195__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08165_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[116\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[108\]
+ net1044 vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout402_A _03566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1144_A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08096_ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[28\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[31\]
+ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[30\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_101_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload80 clknet_leaf_135_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload80/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload91 clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload91/Y sky130_fd_sc_hd__clkinv_4
XANTENNA_fanout1311_A net1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1409_A net1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10206__C net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout771_A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout392_X net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout869_A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08998_ _05303_ _05337_ net603 vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__mux2_4
XANTENNA_fanout657_X net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10960_ _07117_ _07199_ net515 vssd1 vssd1 vccd1 vccd1 _07300_ sky130_fd_sc_hd__mux2_1
XANTENNA__11130__A1 _06920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09874__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11130__B2 _06928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09619_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[24\] net735 _05939_ _05946_
+ _05947_ vssd1 vssd1 vccd1 vccd1 _05959_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout824_X net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10891_ net562 _07208_ _07209_ _07230_ vssd1 vssd1 vccd1 vccd1 _07231_ sky130_fd_sc_hd__a31oi_2
XANTENNA__09730__C net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12630_ net3161 net203 net391 vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_157_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_157_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__14080__B1 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12561_ net3048 net247 net401 vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12864__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14645__A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11621__X _07835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14300_ net1328 vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__inv_2
X_11512_ net1547 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[6\] net877 vssd1 vssd1
+ vccd1 vccd1 _03337_ sky130_fd_sc_hd__mux2_1
XANTENNA__09739__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15280_ net1274 vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12492_ net3097 net219 net409 vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__mux2_1
XANTENNA__08643__A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17729__Q team_01_WB.instance_to_wrap.cpu.f0.write_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_34_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14231_ net1544 vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_117_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13186__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11443_ team_01_WB.instance_to_wrap.cpu.f0.i\[4\] team_01_WB.instance_to_wrap.cpu.f0.i\[3\]
+ _07673_ team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1 _07746_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17528__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14162_ _04188_ _04441_ _04195_ vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__o21a_1
XFILLER_0_34_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11374_ _04478_ _07702_ vssd1 vssd1 vccd1 vccd1 _07703_ sky130_fd_sc_hd__nor2_1
XANTENNA__09177__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10944__A1 _06526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13113_ net1715 net851 net631 team_01_WB.instance_to_wrap.a1.ADR_I\[30\] vssd1 vssd1
+ vccd1 vccd1 _02028_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10325_ net990 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[18\] net951 vssd1
+ vssd1 vccd1 vccd1 _06665_ sky130_fd_sc_hd__and3_1
X_14093_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[5\] _04249_ _04265_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[5\]
+ _04379_ vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__a221o_1
X_13044_ net2465 net2222 net863 vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__mux2_1
X_17921_ net1528 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
XANTENNA__09474__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17678__CLK clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10256_ _06594_ _06595_ vssd1 vssd1 vccd1 vccd1 _06596_ sky130_fd_sc_hd__nand2b_1
Xfanout1210 net1212 vssd1 vssd1 vccd1 vccd1 net1210 sky130_fd_sc_hd__buf_4
Xfanout1221 net1223 vssd1 vssd1 vccd1 vccd1 net1221 sky130_fd_sc_hd__buf_4
X_17852_ clknet_leaf_91_wb_clk_i net1673 _01792_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[122\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1232 net1242 vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12104__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10187_ _06526_ vssd1 vssd1 vccd1 vccd1 _06527_ sky130_fd_sc_hd__inv_2
XANTENNA__10413__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10172__A2 _04636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1243 net1245 vssd1 vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__buf_4
Xfanout1254 net1255 vssd1 vssd1 vccd1 vccd1 net1254 sky130_fd_sc_hd__buf_4
Xfanout1265 net1268 vssd1 vssd1 vccd1 vccd1 net1265 sky130_fd_sc_hd__buf_4
X_16803_ clknet_leaf_26_wb_clk_i _02490_ _00786_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1276 net1277 vssd1 vssd1 vccd1 vccd1 net1276 sky130_fd_sc_hd__buf_4
Xfanout1287 net1289 vssd1 vssd1 vccd1 vccd1 net1287 sky130_fd_sc_hd__buf_4
X_17783_ clknet_leaf_101_wb_clk_i _03459_ _01723_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[53\]
+ sky130_fd_sc_hd__dfstp_1
X_14995_ net1381 vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__inv_2
Xfanout1298 net1301 vssd1 vssd1 vccd1 vccd1 net1298 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11943__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09314__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[22\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16734_ clknet_leaf_85_wb_clk_i _02421_ _00717_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13946_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__or2_2
XFILLER_0_72_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09865__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09640__C net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16665_ clknet_leaf_101_wb_clk_i _02352_ _00648_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11672__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13877_ team_01_WB.EN_VAL_REG net2753 vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__and2b_1
XANTENNA__10880__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15616_ net1233 vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__inv_2
X_12828_ net1851 net641 net609 _03648_ vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14071__B1 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16596_ clknet_leaf_21_wb_clk_i _02283_ _00579_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15547_ net1251 vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__inv_2
XANTENNA__14555__A net1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12759_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] net1060 net363 _03600_
+ vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15478_ net1256 vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__inv_2
XANTENNA__17639__Q team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_17217_ clknet_leaf_54_wb_clk_i _02904_ _01200_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14429_ net1335 vssd1 vssd1 vccd1 vccd1 _00223_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12924__A2 _07752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17148_ clknet_leaf_59_wb_clk_i _02835_ _01131_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_860 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold704 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[15\] vssd1 vssd1 vccd1 vccd1 net2239
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09087__C net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold715 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2250 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold726 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2261 sky130_fd_sc_hd__dlygate4sd3_1
Xhold737 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2272 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_94_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09970_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[3\] net780 net771 _06293_
+ _06298_ vssd1 vssd1 vccd1 vccd1 _06310_ sky130_fd_sc_hd__a2111o_1
Xhold748 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17079_ clknet_leaf_15_wb_clk_i _02766_ _01062_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold759 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2294 sky130_fd_sc_hd__dlygate4sd3_1
X_08921_ net602 _05258_ _05259_ vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_90_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08356__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08852_ net1018 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[3\] net908 vssd1
+ vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__and3_1
XANTENNA__12014__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1404 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2939 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1415 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2950 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10163__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1426 _02149_ vssd1 vssd1 vccd1 vccd1 net2961 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1437 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2972 sky130_fd_sc_hd__dlygate4sd3_1
X_08783_ net1011 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[0\] net882 vssd1
+ vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__and3_1
Xhold1448 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2983 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_140_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1459 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2994 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout185_A net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11853__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09856__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08447__B net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1094_A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10871__A0 _05963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11154__A net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09404_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[27\] net670 net648 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[27\]
+ _05743_ vssd1 vssd1 vccd1 vccd1 _05744_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_9_Left_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14062__B1 _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09335_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[24\] net660 net651 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[24\]
+ _05664_ vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__a221o_1
XANTENNA__12684__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout238_X net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09559__A _05898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09266_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[20\] net671 net646 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08217_ net2945 net2767 net1046 vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__mux2_1
XANTENNA__11601__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09197_ net1004 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[17\] net934 vssd1
+ vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout405_X net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11179__A1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09846__X _06186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08148_ _04583_ _04599_ _04616_ _04617_ vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08044__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09241__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout986_A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08079_ net1768 net570 _04525_ _04553_ vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10110_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[6\] net774 net771 vssd1
+ vssd1 vccd1 vccd1 _06450_ sky130_fd_sc_hd__a21o_1
X_11090_ _04706_ _05835_ _06883_ _07428_ _07429_ vssd1 vssd1 vccd1 vccd1 _07430_ sky130_fd_sc_hd__o311a_1
XFILLER_0_101_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout774_X net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10041_ net994 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[0\] net954 vssd1
+ vssd1 vccd1 vccd1 _06381_ sky130_fd_sc_hd__and3_1
Xhold20 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[4\] vssd1 vssd1 vccd1 vccd1
+ net1555 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10154__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold31 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1566 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[4\] vssd1 vssd1 vccd1 vccd1
+ net1577 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[17\] vssd1 vssd1 vccd1 vccd1
+ net1588 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12859__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout941_X net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold64 _02027_ vssd1 vssd1 vccd1 vccd1 net1599 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13628__B1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold75 _01992_ vssd1 vssd1 vccd1 vccd1 net1610 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11763__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13800_ _01835_ _04176_ _04180_ _04159_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__o22a_1
Xhold86 _01998_ vssd1 vssd1 vccd1 vccd1 net1621 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 net151 vssd1 vssd1 vccd1 vccd1 net1632 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11103__A1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11992_ net575 _07793_ _07951_ vssd1 vssd1 vccd1 vccd1 _07953_ sky130_fd_sc_hd__and3_1
X_14780_ net1249 vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__inv_2
XANTENNA__08638__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13731_ team_01_WB.instance_to_wrap.a1.WRITE_I _04508_ team_01_WB.instance_to_wrap.a1.curr_state\[0\]
+ _04509_ net3089 vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__a32o_1
X_10943_ _07156_ _07282_ net515 vssd1 vssd1 vccd1 vccd1 _07283_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_28_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10862__A0 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16450_ clknet_leaf_52_wb_clk_i _02204_ _00433_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10874_ _05898_ _06779_ _06811_ net512 net548 net537 vssd1 vssd1 vccd1 vccd1 _07214_
+ sky130_fd_sc_hd__mux4_1
X_13662_ net199 net195 _04501_ net645 vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15401_ net1287 vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__inv_2
X_12613_ net2464 net276 net396 vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13593_ _03903_ _04030_ vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12594__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16381_ clknet_leaf_122_wb_clk_i net2610 _00364_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[104\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12544_ net2387 net250 net405 vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15332_ net1221 vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__inv_2
XANTENNA__09469__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08373__A team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09480__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13159__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12475_ net1865 net253 net412 vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__mux2_1
X_15263_ net1314 vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input70_X net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17002_ clknet_leaf_10_wb_clk_i _02689_ _00985_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11426_ _07681_ _07700_ vssd1 vssd1 vccd1 vccd1 _07738_ sky130_fd_sc_hd__nand2_1
XANTENNA__13564__C1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12906__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14214_ net3164 vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_6 _03654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08035__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09232__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15194_ net1370 vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_54_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11938__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14145_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[15\] _04253_ _04258_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[63\]
+ _04429_ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__a221o_1
XANTENNA__10842__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11357_ net1071 _07677_ vssd1 vssd1 vccd1 vccd1 _07686_ sky130_fd_sc_hd__nand2_2
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10393__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10308_ net1129 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[18\] net977
+ vssd1 vssd1 vccd1 vccd1 _06648_ sky130_fd_sc_hd__and3_1
X_14076_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[92\] _04241_ _04267_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[28\]
+ _04363_ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__a221o_1
X_11288_ _04734_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] net1169 vssd1 vssd1
+ vccd1 vccd1 _07628_ sky130_fd_sc_hd__or3b_1
XANTENNA__09635__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17904_ net1439 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
X_13027_ net2538 net2490 net862 vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__mux2_1
X_10239_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[9\] net819 net806 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06579_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_67_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1040 net1041 vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__clkbuf_4
Xfanout1051 net1058 vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__buf_2
X_17835_ clknet_leaf_92_wb_clk_i _03511_ _01775_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[105\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1062 team_01_WB.instance_to_wrap.cpu.RU0.state\[5\] vssd1 vssd1 vccd1 vccd1
+ net1062 sky130_fd_sc_hd__buf_4
Xfanout1073 net1076 vssd1 vssd1 vccd1 vccd1 net1073 sky130_fd_sc_hd__clkbuf_4
Xfanout1084 net1089 vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__buf_1
Xfanout1095 net1096 vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__buf_1
XANTENNA__13454__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17766_ clknet_leaf_99_wb_clk_i _03442_ _01706_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[36\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_107_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14978_ net1346 vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__inv_2
XANTENNA__08548__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16538__Q team_01_WB.instance_to_wrap.cpu.DM0.data_i\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16717_ clknet_leaf_107_wb_clk_i _02404_ _00700_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13929_ _04217_ _04219_ _04220_ vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__and3_4
X_17697_ clknet_leaf_134_wb_clk_i _03381_ _01638_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_77_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16648_ clknet_leaf_62_wb_clk_i _02335_ _00631_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14044__B1 _04266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16579_ clknet_leaf_22_wb_clk_i _02266_ _00562_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_09120_ net1023 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[14\] net924 vssd1
+ vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_44_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09051_ net1029 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[12\] net941 vssd1
+ vssd1 vccd1 vccd1 _05391_ sky130_fd_sc_hd__and3_1
XANTENNA__16273__Q team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08714__C net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12009__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08002_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] vssd1 vssd1 vccd1 vccd1
+ _04500_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold501 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[5\] vssd1 vssd1 vccd1 vccd1
+ net2036 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold512 _02073_ vssd1 vssd1 vccd1 vccd1 net2047 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold523 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2058 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11848__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold534 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2069 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13570__A2 _07251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold545 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2080 sky130_fd_sc_hd__dlygate4sd3_1
Xhold556 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2091 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10384__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold567 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2113 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09953_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[3\] net813 net758 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06293_ sky130_fd_sc_hd__a22o_1
Xhold589 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2124 sky130_fd_sc_hd__dlygate4sd3_1
X_08904_ net1026 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[2\] net924 vssd1
+ vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__and3_1
XANTENNA__12820__X _03643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09884_ net1152 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[5\] net959 vssd1
+ vssd1 vccd1 vccd1 _06224_ sky130_fd_sc_hd__and3_1
XANTENNA__11333__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10136__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1107_A net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1201 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2736 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1212 _03492_ vssd1 vssd1 vccd1 vccd1 net2747 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1223 _02094_ vssd1 vssd1 vccd1 vccd1 net2758 sky130_fd_sc_hd__dlygate4sd3_1
X_08835_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[1\] net689 net659 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__a22o_1
XANTENNA__12679__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1234 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[31\] vssd1 vssd1 vccd1 vccd1
+ net2769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1245 _02105_ vssd1 vssd1 vccd1 vccd1 net2780 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout567_A net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13364__A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1256 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2791 sky130_fd_sc_hd__dlygate4sd3_1
X_08766_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[4\] net699 _05088_ _05092_
+ _05094_ vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__a2111o_1
Xhold1267 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[74\] vssd1 vssd1 vccd1 vccd1
+ net2802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1278 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2813 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09829__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1289 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[103\] vssd1 vssd1 vccd1 vccd1
+ net2824 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08697_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[7\] net699 _05007_ _05025_
+ net708 vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout734_A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1097_X net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10844__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout901_A _04788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09318_ _05657_ vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09289__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10590_ _06897_ _06929_ vssd1 vssd1 vccd1 vccd1 _06930_ sky130_fd_sc_hd__or2_1
XANTENNA__09462__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09249_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[21\] net689 net659 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[21\]
+ _05588_ vssd1 vssd1 vccd1 vccd1 _05589_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_153_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12260_ net2479 net223 net435 vssd1 vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout891_X net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout989_X net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11211_ net530 _07503_ _07549_ net328 vssd1 vssd1 vccd1 vccd1 _07551_ sky130_fd_sc_hd__o211a_1
XANTENNA__08568__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_101_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_142_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13561__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12191_ net2867 net190 net443 vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10515__X _06855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11142_ net375 _06903_ _07014_ _07481_ vssd1 vssd1 vccd1 vccd1 _07482_ sky130_fd_sc_hd__a31o_1
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__buf_2
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__buf_2
X_15950_ net1407 vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__inv_2
X_11073_ _05566_ _06707_ vssd1 vssd1 vccd1 vccd1 _07413_ sky130_fd_sc_hd__or2_1
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 ADR_O[30] sky130_fd_sc_hd__buf_2
X_10024_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[1\] net778 _06362_ _06363_
+ vssd1 vssd1 vccd1 vccd1 _06364_ sky130_fd_sc_hd__a211o_1
X_14901_ net1275 vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__inv_2
XANTENNA_input30_A DAT_I[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12589__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15881_ net1347 vssd1 vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_129_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17620_ clknet_leaf_2_wb_clk_i _03305_ _01561_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10250__X _06590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14832_ net1250 vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__inv_2
XANTENNA__14089__B net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_17 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17551_ clknet_leaf_34_wb_clk_i _03238_ _01534_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_101_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_101_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12824__A1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14763_ net1346 vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__inv_2
X_11975_ net2104 net263 net472 vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__mux2_1
XANTENNA__12824__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16502_ clknet_leaf_2_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[0\]
+ _00485_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13714_ _04102_ _04119_ _04126_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[5\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10926_ _06980_ _07227_ vssd1 vssd1 vccd1 vccd1 _07266_ sky130_fd_sc_hd__nor2_1
X_17482_ clknet_leaf_9_wb_clk_i _03169_ _01465_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14026__B1 _04258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14694_ net1195 vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__inv_2
X_16433_ clknet_leaf_141_wb_clk_i _02187_ _00416_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10857_ net370 _07195_ _07196_ net340 _04970_ vssd1 vssd1 vccd1 vccd1 _07197_ sky130_fd_sc_hd__o32a_1
X_13645_ net989 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] _04079_ _04080_
+ vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08815__B net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_140_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16364_ clknet_leaf_97_wb_clk_i _02118_ _00347_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[87\]
+ sky130_fd_sc_hd__dfrtp_1
X_10788_ net335 _07127_ _07126_ vssd1 vssd1 vccd1 vccd1 _07128_ sky130_fd_sc_hd__o21ai_1
X_13576_ net724 _07231_ net986 vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09453__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15315_ net1392 vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__inv_2
X_12527_ net2810 net212 net404 vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__mux2_1
XANTENNA__15929__A net1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16295_ clknet_leaf_101_wb_clk_i _02049_ _00278_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_15246_ net1297 vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08831__A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12458_ net2085 net224 net411 vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08559__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11409_ _07701_ _07711_ _07727_ net323 vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15177_ net1293 vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__inv_2
X_12389_ net3141 net288 net424 vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12760__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14128_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[86\] _04245_ _04396_ _04152_
+ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__a211o_1
XFILLER_0_123_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14059_ _04347_ vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__inv_2
XANTENNA__10118__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12499__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08620_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[11\] net665 net654 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[11\]
+ _04959_ vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__a221o_1
XANTENNA__08731__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17818_ clknet_leaf_122_wb_clk_i net2877 _01758_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[88\]
+ sky130_fd_sc_hd__dfrtp_1
X_08551_ net1077 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[19\] net891
+ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__and3_1
XANTENNA__08709__C net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17749_ clknet_leaf_96_wb_clk_i _03425_ _01689_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10826__A0 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08482_ net1004 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[23\] net882 vssd1
+ vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09692__B1 _06030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10841__A3 _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_99_Left_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09103_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[13\] net688 _05431_
+ _05433_ _05440_ vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08444__C net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12962__S net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12815__X _03639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_131_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1057_A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13528__C1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09034_ _05339_ _05373_ net603 vssd1 vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__mux2_4
XANTENNA__08741__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13543__A2 _07111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold320 team_01_WB.instance_to_wrap.cpu.f0.write_data\[23\] vssd1 vssd1 vccd1 vccd1
+ net1855 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold331 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1866 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08460__B net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold342 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1877 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1224_A net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold353 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[127\] vssd1 vssd1 vccd1 vccd1
+ net1888 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 net139 vssd1 vssd1 vccd1 vccd1 net1899 sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1910 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold386 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1921 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout800 net801 vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout684_A _04780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold397 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1932 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout811 net814 vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__clkbuf_8
X_09936_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[4\] net812 net798 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[4\]
+ _06275_ vssd1 vssd1 vccd1 vccd1 _06276_ sky130_fd_sc_hd__a221o_1
Xfanout822 net824 vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10109__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11306__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout833 net834 vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__buf_1
Xfanout844 net845 vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__buf_2
Xfanout855 net858 vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__clkbuf_4
Xfanout866 net867 vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__clkbuf_2
X_09867_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[12\] net741 _06205_ _06206_
+ vssd1 vssd1 vccd1 vccd1 _06207_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout472_X net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout877 team_01_WB.instance_to_wrap.cpu.DM0.next_enable vssd1 vssd1 vccd1 vccd1
+ net877 sky130_fd_sc_hd__clkbuf_4
Xfanout888 _04799_ vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__buf_2
Xhold1020 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2555 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout899 _04793_ vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__buf_2
Xhold1031 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2566 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout949_A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1042 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2577 sky130_fd_sc_hd__dlygate4sd3_1
X_08818_ net1105 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[1\] net880 vssd1
+ vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__and3_1
XANTENNA__12202__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1053 _03433_ vssd1 vssd1 vccd1 vccd1 net2588 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09798_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[14\] net789 net740 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06138_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_107_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1064 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2599 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1075 _02135_ vssd1 vssd1 vccd1 vccd1 net2610 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1086 _02053_ vssd1 vssd1 vccd1 vccd1 net2621 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1097 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2632 sky130_fd_sc_hd__dlygate4sd3_1
X_08749_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[4\] net932 vssd1
+ vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout737_X net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12806__B2 _03632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10817__A0 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ net2112 net223 net495 vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__mux2_1
XANTENNA__08475__X _04815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14008__B1 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09683__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10711_ net557 _07050_ vssd1 vssd1 vccd1 vccd1 _07051_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_155_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout904_X net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11691_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] _07805_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\]
+ vssd1 vssd1 vccd1 vccd1 _07890_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_120_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11342__A team_01_WB.instance_to_wrap.cpu.f0.i\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10642_ _06129_ net371 net549 vssd1 vssd1 vccd1 vccd1 _06982_ sky130_fd_sc_hd__mux2_1
X_13430_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] net595 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\]
+ vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09435__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13361_ _04484_ _07683_ vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_3_5_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12872__S net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10573_ _04741_ _04743_ vssd1 vssd1 vccd1 vccd1 _06913_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15100_ net1244 vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__inv_2
X_12312_ net2843 net228 net431 vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__mux2_1
X_13292_ team_01_WB.instance_to_wrap.cpu.f0.i\[23\] _03744_ vssd1 vssd1 vccd1 vccd1
+ _03778_ sky130_fd_sc_hd__nand2_1
X_16080_ clknet_leaf_130_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[2\]
+ _00068_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__08651__A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17737__Q team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12243_ net2634 net258 net441 vssd1 vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__mux2_1
X_15031_ net1220 vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__inv_2
XANTENNA__08370__B team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12742__B1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12174_ net2327 net230 net449 vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__mux2_1
XANTENNA__09185__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11125_ net535 _07453_ vssd1 vssd1 vccd1 vccd1 _07465_ sky130_fd_sc_hd__nand2_1
XANTENNA__08961__A2 _05300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16982_ clknet_leaf_30_wb_clk_i _02669_ _00965_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_15933_ net1417 vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__inv_2
X_11056_ net555 _06280_ vssd1 vssd1 vccd1 vccd1 _07396_ sky130_fd_sc_hd__nand2_1
XANTENNA__09910__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10007_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[1\] net820 net812 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06347_ sky130_fd_sc_hd__a22o_1
X_15864_ net1347 vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__inv_2
XANTENNA__12112__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10520__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17603_ clknet_leaf_86_wb_clk_i _03290_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_14815_ net1317 vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__inv_2
XANTENNA__08529__C net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15795_ net1231 vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11951__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14828__A net1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17534_ clknet_leaf_79_wb_clk_i _03221_ _01517_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14746_ net1189 vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__inv_2
X_11958_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\] team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\]
+ vssd1 vssd1 vccd1 vccd1 _07951_ sky130_fd_sc_hd__and2b_2
XANTENNA__08826__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17465_ clknet_leaf_103_wb_clk_i _03152_ _01448_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10909_ _07100_ _07242_ _07248_ net327 _07247_ vssd1 vssd1 vccd1 vccd1 _07249_ sky130_fd_sc_hd__a221o_1
X_14677_ net1227 vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__inv_2
X_11889_ net1928 net317 net486 vssd1 vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16416_ clknet_leaf_124_wb_clk_i _02170_ _00399_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13628_ net722 _07269_ net1074 vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__o21a_1
XFILLER_0_7_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17396_ clknet_leaf_22_wb_clk_i _03083_ _01379_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09426__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13222__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_55_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15659__A net1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16347_ clknet_leaf_118_wb_clk_i net2919 _00330_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[70\]
+ sky130_fd_sc_hd__dfrtp_1
X_13559_ net185 _04007_ _04008_ net723 vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__a211o_1
XFILLER_0_14_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14563__A net1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10587__A2 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09657__A net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16278_ clknet_leaf_123_wb_clk_i _02032_ _00261_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08561__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10992__C1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18017_ net637 vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13525__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15229_ net1311 vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10155__X _06495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11536__B2 net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09095__C net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08952__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15394__A net1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07982_ team_01_WB.instance_to_wrap.cpu.f0.i\[14\] vssd1 vssd1 vccd1 vccd1 _04480_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_10_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10034__C net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09721_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[21\] net757 _06043_ _06044_
+ _06046_ vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_129_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12022__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09652_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[23\] net782 _05970_ _05971_
+ _05977_ vssd1 vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10511__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08603_ _04935_ _04936_ _04939_ _04942_ vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__or4_2
X_09583_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[25\] net822 net751 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11861__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08534_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[18\] net648 _04848_
+ _04851_ _04857_ vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13997__C1 net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10985__B _06398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11472__B1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08465_ net1083 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[23\] net883
+ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout432_A _07964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1174_A team_01_WB.instance_to_wrap.cpu.DM0.ihit vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08396_ _04733_ _04735_ _04734_ _04731_ vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_147_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout220_X net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12692__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09567__A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09017_ net1012 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[9\] net878 vssd1
+ vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout899_A _04793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08902__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13516__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11527__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold150 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1685 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold161 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1
+ net1696 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10735__C1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold172 _01987_ vssd1 vssd1 vccd1 vccd1 net1707 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout687_X net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold183 _02024_ vssd1 vssd1 vccd1 vccd1 net1718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 team_01_WB.instance_to_wrap.a1.ADR_I\[14\] vssd1 vssd1 vccd1 vccd1 net1729
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout630 _03738_ vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__buf_2
Xfanout641 _03572_ vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__clkbuf_2
X_09919_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[4\] net785 net760 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06259_ sky130_fd_sc_hd__a22o_1
Xfanout652 _04819_ vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__buf_6
Xfanout663 _04806_ vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__clkbuf_8
Xfanout674 _04791_ vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__buf_6
Xfanout685 _04780_ vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_126_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12930_ net356 _03695_ _03696_ net869 net2467 vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__a32o_1
Xfanout696 _04766_ vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10502__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08349__C net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11056__B _06280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12861_ net2313 net311 net380 vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_923 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11771__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14600_ net1356 vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_1_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ net2260 net227 net491 vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__mux2_1
X_15580_ net1248 vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__inv_2
XANTENNA__08646__A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09656__B1 _05994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12792_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[12\] _07520_ net1034 vssd1 vssd1
+ vccd1 vccd1 _03623_ sky130_fd_sc_hd__mux2_1
X_14531_ net1417 vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__inv_2
X_11743_ net716 net321 vssd1 vssd1 vccd1 vccd1 _07932_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17250_ clknet_leaf_58_wb_clk_i _02937_ _01233_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_14462_ net1225 vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09408__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11674_ _07874_ _07876_ net611 vssd1 vssd1 vccd1 vccd1 _07877_ sky130_fd_sc_hd__mux2_2
XFILLER_0_83_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16201_ clknet_leaf_159_wb_clk_i _01961_ _00189_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13413_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] _05116_ _07641_ _07640_
+ vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__a31o_1
X_17181_ clknet_leaf_64_wb_clk_i _02868_ _01164_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10625_ net528 net503 vssd1 vssd1 vccd1 vccd1 _06965_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14393_ net1186 vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16132_ clknet_leaf_127_wb_clk_i _00023_ _00120_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.state\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__12963__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13344_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[15\] net827 _03816_ _03818_
+ vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__o22a_1
X_10556_ net545 _05899_ _06895_ vssd1 vssd1 vccd1 vccd1 _06896_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10974__C1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16063_ clknet_leaf_3_wb_clk_i _01856_ _00051_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_45_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12107__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13275_ net587 _03763_ _03764_ net564 vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__a22o_1
X_10487_ _05869_ _05870_ vssd1 vssd1 vccd1 vccd1 _06827_ sky130_fd_sc_hd__or2_1
XANTENNA__10416__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11518__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15014_ net1381 vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__inv_2
X_12226_ net3113 net190 net439 vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__mux2_1
XANTENNA__11946__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12157_ _07791_ net576 _07942_ vssd1 vssd1 vccd1 vccd1 _07958_ sky130_fd_sc_hd__and3_4
XANTENNA__12190__X _07959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11108_ _07071_ _07447_ _07444_ _07441_ vssd1 vssd1 vccd1 vccd1 _07448_ sky130_fd_sc_hd__o211a_1
X_12088_ net2287 net319 net462 vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__mux2_1
X_16965_ clknet_leaf_51_wb_clk_i _02652_ _00948_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11039_ _07259_ _07373_ _07377_ _07378_ vssd1 vssd1 vccd1 vccd1 _07379_ sky130_fd_sc_hd__and4b_1
X_15916_ net1360 vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__inv_2
X_16896_ clknet_leaf_39_wb_clk_i _02583_ _00879_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09895__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15847_ net1326 vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15778_ net1197 vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__inv_2
XANTENNA__09647__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08556__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09151__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09111__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17517_ clknet_leaf_68_wb_clk_i _03204_ _01500_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14729_ net1209 vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08250_ net2714 net2591 net1047 vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__mux2_1
X_17448_ clknet_leaf_63_wb_clk_i _03135_ _01431_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08181_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[100\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[92\]
+ net1044 vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17379_ clknet_leaf_26_wb_clk_i _03066_ _01362_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_9_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_31_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08722__C net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12017__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10326__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09178__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_151_Right_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11856__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09704_ net1154 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[21\] net959
+ vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_143_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09350__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09635_ net1135 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[23\] net948
+ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout647_A _04825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09566_ net1149 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[25\] net974
+ vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11604__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08517_ net1079 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[18\] net922
+ vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__and3_1
XFILLER_0_148_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13985__A2 _04226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09497_ _04706_ _05836_ vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout435_X net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1177_X net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11323__C team_01_WB.instance_to_wrap.cpu.DM0.data_i\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08448_ net1121 net1124 net1127 net1118 vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__and4b_4
XFILLER_0_93_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13198__B1 _03738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15299__A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08379_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[4\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\]
+ net1170 vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__and3b_1
XANTENNA_fanout602_X net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1344_X net1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11748__A1 _07489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10410_ _06748_ _06749_ _05934_ _05967_ vssd1 vssd1 vccd1 vccd1 _06750_ sky130_fd_sc_hd__a211o_2
XANTENNA__09297__A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11390_ _07717_ _07718_ _04465_ vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09810__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08632__C net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10341_ net991 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[17\] net962 vssd1
+ vssd1 vccd1 vccd1 _06681_ sky130_fd_sc_hd__and3_1
XFILLER_0_143_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09169__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13060_ net2569 net2046 net864 vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__mux2_1
X_10272_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[19\] net739 _06609_ _06610_
+ _06611_ vssd1 vssd1 vccd1 vccd1 _06612_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_143_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout971_X net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12011_ net2607 net253 net467 vssd1 vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__mux2_1
XANTENNA__11766__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08916__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13855__A_N net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13370__B1 _07650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1403 net1409 vssd1 vssd1 vccd1 vccd1 net1403 sky130_fd_sc_hd__buf_2
Xfanout1414 net1428 vssd1 vssd1 vccd1 vccd1 net1414 sky130_fd_sc_hd__buf_2
Xfanout1425 net1428 vssd1 vssd1 vccd1 vccd1 net1425 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout460 _07955_ vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout471 _07952_ vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__buf_6
Xfanout482 _07949_ vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__clkbuf_4
X_16750_ clknet_leaf_27_wb_clk_i _02437_ _00733_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13962_ _04218_ _04242_ vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__nor2_4
Xfanout493 _07944_ vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13673__A1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11133__C1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13673__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15701_ net1293 vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_79_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09341__A2 _05678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12913_ _04881_ net578 vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__nor2_1
X_16681_ clknet_leaf_35_wb_clk_i _02368_ _00664_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12597__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13893_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[0\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[1\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[2\] vssd1 vssd1 vccd1 vccd1 _04198_
+ sky130_fd_sc_hd__a21o_1
X_15632_ net1251 vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__inv_2
X_12844_ net2823 net241 net380 vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__mux2_1
XANTENNA__08807__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15563_ net1424 vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12775_ net1722 net638 net606 _03611_ vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17302_ clknet_leaf_24_wb_clk_i _02989_ _01285_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14514_ net1363 vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11726_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[6\] net716 vssd1 vssd1 vccd1
+ vccd1 _07918_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15494_ net1380 vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13189__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17233_ clknet_leaf_112_wb_clk_i _02920_ _01216_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_14445_ net1225 vssd1 vssd1 vccd1 vccd1 _00239_ sky130_fd_sc_hd__inv_2
X_11657_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[20\] net713 vssd1 vssd1 vccd1
+ vccd1 _07863_ sky130_fd_sc_hd__or2_1
XANTENNA__11739__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10608_ _06946_ _06947_ vssd1 vssd1 vccd1 vccd1 _06948_ sky130_fd_sc_hd__nor2_1
X_17164_ clknet_leaf_147_wb_clk_i _02851_ _01147_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_14376_ net1208 vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__inv_2
XANTENNA__09638__C net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11588_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] _07803_ vssd1 vssd1
+ vccd1 vccd1 _07805_ sky130_fd_sc_hd__and2_1
XFILLER_0_101_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16115_ clknet_leaf_136_wb_clk_i _01890_ _00103_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_52_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold908 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2443 sky130_fd_sc_hd__dlygate4sd3_1
X_13327_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[19\] net826 _03805_ vssd1 vssd1
+ vccd1 vccd1 _01887_ sky130_fd_sc_hd__o21a_1
X_10539_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[31\] net688 net670 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06879_ sky130_fd_sc_hd__a22o_1
Xhold919 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[118\] vssd1 vssd1 vccd1 vccd1
+ net2454 sky130_fd_sc_hd__dlygate4sd3_1
X_17095_ clknet_leaf_106_wb_clk_i _02782_ _01078_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16046_ clknet_leaf_158_wb_clk_i _01839_ _00034_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.BUSY_O
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13258_ team_01_WB.instance_to_wrap.cpu.f0.i\[28\] _03749_ vssd1 vssd1 vccd1 vccd1
+ _03750_ sky130_fd_sc_hd__nand2_1
XANTENNA__11676__S net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12209_ net1903 net253 net443 vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10175__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13189_ net20 net837 net630 net2115 vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__a22o_1
XANTENNA__11911__A1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11248__Y _07588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09580__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17997_ net1506 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__buf_2
Xhold1608 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net3143 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1619 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net3154 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13113__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16948_ clknet_leaf_22_wb_clk_i _02635_ _00931_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13664__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16879_ clknet_leaf_35_wb_clk_i _02566_ _00862_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_09420_ net559 _05759_ _05737_ vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__o21ai_2
XANTENNA__12300__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08717__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11427__B1 _07699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09351_ _05689_ _05690_ vssd1 vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__or2_1
XANTENNA__11978__A1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08302_ net1144 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[30\] net972
+ vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09282_ net1084 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[22\] net939
+ vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08233_ net2616 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[40\] net1049 vssd1 vssd1
+ vccd1 vccd1 _03454_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10650__A1 _06811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_99_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout228_A _07900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09399__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08164_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[117\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[109\]
+ net1051 vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08452__C net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08095_ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[25\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[24\]
+ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[27\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__or4_1
XANTENNA__12823__X _03645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload70 clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload70/Y sky130_fd_sc_hd__clkinv_8
XANTENNA_fanout1137_A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload81 clknet_leaf_136_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload81/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__14144__A2 _04244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload92 clknet_leaf_143_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload92/Y sky130_fd_sc_hd__inv_6
XFILLER_0_140_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout597_A net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10166__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1304_A net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09283__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08997_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[8\] net702 _05320_ _05336_
+ vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__a2bb2o_4
XANTENNA_fanout764_A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout385_X net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09859__B1 _04678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13655__A1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09323__A2 _04766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout931_A net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13814__B net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11615__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09618_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[24\] net795 net775 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__a22o_1
XANTENNA__12210__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10890_ _07054_ _07228_ _07229_ vssd1 vssd1 vccd1 vccd1 _07230_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09549_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[28\] net800 net773 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[28\]
+ _05884_ vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__a221o_1
XANTENNA__11969__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout817_X net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11053__C net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12560_ net2470 net210 net399 vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__mux2_1
XANTENNA__08483__X _04823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11511_ net1699 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[7\] net876 vssd1 vssd1
+ vccd1 vccd1 _03338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12491_ net1704 net224 net407 vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__mux2_1
XANTENNA__12918__B1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14230_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[2\] vssd1 vssd1 vccd1
+ vccd1 _02257_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11442_ _07676_ _07745_ vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_126_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_126_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_22_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11197__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08598__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13591__B1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14161_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[3\] _04187_ vssd1 vssd1 vccd1
+ vccd1 _04441_ sky130_fd_sc_hd__nor2_1
X_11373_ team_01_WB.instance_to_wrap.cpu.f0.i\[15\] _07682_ vssd1 vssd1 vccd1 vccd1
+ _07702_ sky130_fd_sc_hd__nand2_1
XANTENNA__12733__X _03583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10944__A2 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input60_A wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13112_ net1774 net843 net631 team_01_WB.instance_to_wrap.a1.ADR_I\[31\] vssd1 vssd1
+ vccd1 vccd1 _02029_ sky130_fd_sc_hd__a22o_1
X_10324_ net1135 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[18\] net963
+ vssd1 vssd1 vccd1 vccd1 _06664_ sky130_fd_sc_hd__and3_1
XANTENNA__14135__A2 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14092_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[29\] _04267_ _04268_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[77\]
+ vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__a22o_1
XANTENNA__13277__A team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17920_ net1527 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
X_10255_ net339 _06593_ vssd1 vssd1 vccd1 vccd1 _06595_ sky130_fd_sc_hd__nand2_1
X_13043_ net2541 net2480 net861 vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_57_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1200 net1201 vssd1 vssd1 vccd1 vccd1 net1200 sky130_fd_sc_hd__buf_2
Xfanout1211 net1212 vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__buf_2
X_17851_ clknet_leaf_93_wb_clk_i net1650 _01791_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09193__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11509__B _07756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10186_ net626 _06525_ _06502_ vssd1 vssd1 vccd1 vccd1 _06526_ sky130_fd_sc_hd__o21ai_4
Xfanout1222 net1223 vssd1 vssd1 vccd1 vccd1 net1222 sky130_fd_sc_hd__buf_2
Xfanout1233 net1235 vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1244 net1245 vssd1 vssd1 vccd1 vccd1 net1244 sky130_fd_sc_hd__buf_4
X_16802_ clknet_leaf_57_wb_clk_i _02489_ _00785_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1255 net1303 vssd1 vssd1 vccd1 vccd1 net1255 sky130_fd_sc_hd__clkbuf_4
Xfanout1266 net1268 vssd1 vssd1 vccd1 vccd1 net1266 sky130_fd_sc_hd__buf_4
X_17782_ clknet_leaf_99_wb_clk_i _03458_ _01722_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[52\]
+ sky130_fd_sc_hd__dfstp_1
X_14994_ net1290 vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__inv_2
Xfanout1277 net1302 vssd1 vssd1 vccd1 vccd1 net1277 sky130_fd_sc_hd__buf_2
Xfanout1288 net1289 vssd1 vssd1 vccd1 vccd1 net1288 sky130_fd_sc_hd__buf_4
Xfanout290 net291 vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__clkbuf_2
Xfanout1299 net1301 vssd1 vssd1 vccd1 vccd1 net1299 sky130_fd_sc_hd__buf_4
XANTENNA__09314__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16733_ clknet_leaf_69_wb_clk_i _02420_ _00716_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13945_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__nor2_2
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12120__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16664_ clknet_leaf_38_wb_clk_i _02351_ _00647_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13876_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[13\] _04186_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[14\]
+ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.lcd_en sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15615_ net1311 vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__inv_2
XANTENNA__10880__A1 _05566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09078__A1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12827_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] net1063 net365 _03647_
+ vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__a22o_1
X_16595_ clknet_leaf_149_wb_clk_i _02282_ _00578_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15546_ net1370 vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12758_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[23\] _07111_ net1034 vssd1 vssd1
+ vccd1 vccd1 _03600_ sky130_fd_sc_hd__mux2_1
XANTENNA__08834__A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11709_ net2029 net251 net500 vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15477_ net1282 vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_62_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12689_ net1926 net223 net383 vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17216_ clknet_leaf_48_wb_clk_i _02903_ _01199_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12909__B1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14428_ net1305 vssd1 vssd1 vccd1 vccd1 _00222_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08589__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_96_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17147_ clknet_leaf_74_wb_clk_i _02834_ _01130_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13582__B1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold705 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2240 sky130_fd_sc_hd__dlygate4sd3_1
X_14359_ net1326 vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__inv_2
XANTENNA__14571__A net1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold716 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2251 sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2262 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10307__C net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold738 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2273 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14126__A2 _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold749 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2284 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17078_ clknet_leaf_12_wb_clk_i _02765_ _01061_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16029_ net1309 vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__inv_2
X_08920_ net602 _05258_ _05259_ vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__a21o_1
XANTENNA__10148__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08851_ net1098 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[3\] net912 vssd1
+ vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_71_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1405 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2940 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1416 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2951 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1427 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2962 sky130_fd_sc_hd__dlygate4sd3_1
X_08782_ net1011 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[0\] net896 vssd1
+ vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__and3_1
Xhold1438 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2973 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10042__C net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1449 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2984 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_140_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09305__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12030__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09403_ net1080 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[27\] net906
+ net664 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[27\] vssd1 vssd1 vccd1
+ vccd1 _05743_ sky130_fd_sc_hd__a32o_1
XANTENNA__10871__A1 _05996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout345_A net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1087_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09334_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[24\] net694 _05673_
+ net706 vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__a211o_1
XANTENNA__08744__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_80_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09265_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[20\] _04778_ net685 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[20\]
+ _05597_ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__a221o_1
X_08216_ net2675 net2529 net1056 vssd1 vssd1 vccd1 vccd1 _03471_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09196_ net1005 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[17\] net896 vssd1
+ vssd1 vccd1 vccd1 _05536_ sky130_fd_sc_hd__and3_1
XFILLER_0_43_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08147_ _04465_ team_01_WB.instance_to_wrap.cpu.f0.num\[31\] team_01_WB.instance_to_wrap.cpu.f0.num\[25\]
+ _04470_ _04585_ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__o221a_1
XANTENNA__10387__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08044__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08078_ team_01_WB.instance_to_wrap.cpu.f0.i\[3\] team_01_WB.instance_to_wrap.cpu.K0.keyvalid
+ _04523_ _04552_ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__a31o_1
XANTENNA__14117__A2 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13809__B net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout881_A _04810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13097__A net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout979_A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12205__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10139__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10040_ net1142 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[0\] net968 vssd1
+ vssd1 vccd1 vccd1 _06380_ sky130_fd_sc_hd__and3_1
XANTENNA__09544__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold10 team_01_WB.instance_to_wrap.a1.ADR_I\[17\] vssd1 vssd1 vccd1 vccd1 net1545
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout767_X net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold21 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1556 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[7\] vssd1 vssd1 vccd1 vccd1 net1567
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13628__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold43 team_01_WB.instance_to_wrap.cpu.f0.write_data\[1\] vssd1 vssd1 vccd1 vccd1
+ net1578 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[24\] vssd1 vssd1 vccd1 vccd1 net1589
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 team_01_WB.instance_to_wrap.cpu.f0.write_data\[13\] vssd1 vssd1 vccd1 vccd1
+ net1600 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08919__A net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold76 net118 vssd1 vssd1 vccd1 vccd1 net1611 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11639__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11616__Y _07831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold87 net104 vssd1 vssd1 vccd1 vccd1 net1622 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout934_X net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11991_ net2154 net288 net472 vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__mux2_1
Xhold98 team_01_WB.instance_to_wrap.cpu.f0.write_data\[9\] vssd1 vssd1 vccd1 vccd1
+ net1633 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09741__C net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11103__A2 _06280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11345__A team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_98_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13730_ team_01_WB.instance_to_wrap.cpu.DM0.state\[0\] _04132_ _04133_ net1175 vssd1
+ vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__a22o_1
X_10942_ _06636_ _06671_ _06707_ _06738_ net549 net538 vssd1 vssd1 vccd1 vccd1 _07282_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10311__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11064__B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_119_Left_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13661_ _03874_ _03875_ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__xor2_1
XFILLER_0_151_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12875__S net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10873_ net530 _07212_ vssd1 vssd1 vccd1 vccd1 _07213_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14656__A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15400_ net1376 vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12612_ net2099 net303 net396 vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16380_ clknet_leaf_96_wb_clk_i _02134_ _00363_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[103\]
+ sky130_fd_sc_hd__dfrtp_1
X_13592_ net987 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] _04035_ _04036_
+ vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_130_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08654__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15331_ net1250 vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12543_ net2589 net227 net403 vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__mux2_1
XANTENNA__08373__B team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15262_ net1345 vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__inv_2
X_12474_ net2751 net258 net414 vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17001_ clknet_leaf_38_wb_clk_i _02688_ _00984_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17645__CLK clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14213_ net2574 vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__clkbuf_1
X_11425_ team_01_WB.instance_to_wrap.cpu.f0.i\[9\] _07736_ vssd1 vssd1 vccd1 vccd1
+ _07737_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15193_ net1238 vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__inv_2
XANTENNA__10378__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_7 _03654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14144_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[103\] _04244_ _04245_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[87\]
+ vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_128_Left_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11356_ _04483_ _07684_ vssd1 vssd1 vccd1 vccd1 _07685_ sky130_fd_sc_hd__nor2_1
XANTENNA__09783__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10307_ net1129 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[18\] net956
+ vssd1 vssd1 vccd1 vccd1 _06647_ sky130_fd_sc_hd__and3_1
XANTENNA__12115__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14075_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[44\] _04246_ _04252_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[108\]
+ vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__a22o_1
X_11287_ _06961_ _07622_ _07625_ _07626_ vssd1 vssd1 vccd1 vccd1 _07627_ sky130_fd_sc_hd__or4_2
XFILLER_0_120_886 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_94_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13026_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[60\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[68\]
+ net855 vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__mux2_1
X_17903_ net1438 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
X_10238_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[9\] net781 net772 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06578_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_4_0__f_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1030 net1031 vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11954__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1041 team_01_WB.instance_to_wrap.cpu.RU0.InstrRead vssd1 vssd1 vccd1 vccd1
+ net1041 sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_23_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10169_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[10\] _04654_ net750
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[10\] vssd1 vssd1 vccd1 vccd1
+ _06509_ sky130_fd_sc_hd__a22o_1
Xfanout1052 net1058 vssd1 vssd1 vccd1 vccd1 net1052 sky130_fd_sc_hd__clkbuf_4
X_17834_ clknet_leaf_122_wb_clk_i _03510_ _01774_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[104\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1063 team_01_WB.instance_to_wrap.cpu.RU0.state\[5\] vssd1 vssd1 vccd1 vccd1
+ net1063 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08829__A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1074 net1076 vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_156_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1085 net1088 vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__clkbuf_2
Xfanout1096 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[24\] vssd1 vssd1 vccd1 vccd1
+ net1096 sky130_fd_sc_hd__buf_2
X_14977_ net1280 vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__inv_2
X_17765_ clknet_leaf_97_wb_clk_i _03441_ _01705_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13928_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__and2_2
X_16716_ clknet_leaf_19_wb_clk_i _02403_ _00699_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_137_Left_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17696_ clknet_leaf_134_wb_clk_i _03380_ _01637_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10302__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16647_ clknet_leaf_99_wb_clk_i _02334_ _00630_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13859_ net1177 net1064 net3184 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[20\]
+ sky130_fd_sc_hd__and3b_1
XANTENNA__13470__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16578_ clknet_leaf_75_wb_clk_i _02265_ _00561_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15529_ net1295 vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09050_ net1109 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[12\] net912
+ vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__and3_1
XANTENNA__10081__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09098__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08001_ net1073 vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12814__A net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold502 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2037 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10037__C net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold513 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2048 sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2059 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09774__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold535 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2070 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09826__C net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold546 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2081 sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2092 sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[11\] vssd1 vssd1 vccd1 vccd1
+ net2103 sky130_fd_sc_hd__dlygate4sd3_1
X_09952_ net1154 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[3\] net982 vssd1
+ vssd1 vccd1 vccd1 _06292_ sky130_fd_sc_hd__and3_1
Xhold579 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2114 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11318__C1 _07650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08903_ net1026 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[2\] net936 vssd1
+ vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__and3_1
XANTENNA__09526__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09883_ net1153 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[5\] net969 vssd1
+ vssd1 vccd1 vccd1 _06223_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout295_A _07926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11864__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08734__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1202 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[54\] vssd1 vssd1 vccd1 vccd1
+ net2737 sky130_fd_sc_hd__dlygate4sd3_1
X_08834_ net1022 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[1\] net884 vssd1
+ vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1213 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2748 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08739__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1224 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2759 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1002_A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1235 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2770 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1246 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1257 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2792 sky130_fd_sc_hd__dlygate4sd3_1
X_08765_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[4\] net678 _05078_ _05096_
+ net707 vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__a2111o_1
Xhold1268 _02113_ vssd1 vssd1 vccd1 vccd1 net2803 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout462_A _07955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1279 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2814 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08696_ _05032_ _05033_ _05034_ _05035_ vssd1 vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__or4_2
XANTENNA__10500__C net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10844__A1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12695__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout727_A net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08474__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08905__C net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09317_ net597 _05654_ _05656_ vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__o21a_2
XANTENNA_fanout515_X net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09248_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[21\] net675 net673 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09179_ net1010 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[16\] net896 vssd1
+ vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__and3_1
XANTENNA__10943__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11210_ net338 _07043_ _07548_ net557 vssd1 vssd1 vccd1 vccd1 _07550_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12190_ _07790_ _07791_ net575 vssd1 vssd1 vccd1 vccd1 _07959_ sky130_fd_sc_hd__and3_4
XANTENNA_fanout884_X net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09736__C net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08640__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11141_ net370 _07479_ _07480_ _07389_ vssd1 vssd1 vccd1 vccd1 _07481_ sky130_fd_sc_hd__o31a_1
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__buf_2
X_11072_ _07403_ _07406_ _07407_ _07411_ _07364_ vssd1 vssd1 vccd1 vccd1 _07412_ sky130_fd_sc_hd__a41o_1
XANTENNA__09517__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__buf_2
XANTENNA__12730__Y _03580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 ADR_O[31] sky130_fd_sc_hd__buf_2
XANTENNA__11774__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10023_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[1\] net816 net805 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06363_ sky130_fd_sc_hd__a22o_1
X_14900_ net1378 vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__inv_2
X_15880_ net1349 vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__inv_2
XANTENNA__10532__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08649__A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17922__1529 vssd1 vssd1 vccd1 vccd1 net1529 _17922__1529/LO sky130_fd_sc_hd__conb_1
XFILLER_0_99_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14831_ net1299 vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__inv_2
XANTENNA_input23_A DAT_I[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09471__C net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17550_ clknet_leaf_28_wb_clk_i _03237_ _01533_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_14762_ net1370 vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__inv_2
X_11974_ net1780 net265 net471 vssd1 vssd1 vccd1 vccd1 _03008_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16501_ clknet_leaf_157_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_read_i
+ _00484_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.READ_I sky130_fd_sc_hd__dfrtp_1
X_13713_ team_01_WB.instance_to_wrap.cpu.c0.count\[4\] _04101_ team_01_WB.instance_to_wrap.cpu.c0.count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__a21o_1
X_17481_ clknet_leaf_35_wb_clk_i _03168_ _01464_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10925_ net524 _07215_ vssd1 vssd1 vccd1 vccd1 _07265_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14693_ net1198 vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__inv_2
X_16432_ clknet_leaf_135_wb_clk_i _02186_ _00415_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_141_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_141_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13644_ net722 _07323_ net1075 vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__o21a_1
X_10856_ net337 _06918_ _07194_ vssd1 vssd1 vccd1 vccd1 _07196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16363_ clknet_leaf_119_wb_clk_i _02117_ _00346_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[86\]
+ sky130_fd_sc_hd__dfrtp_1
X_13575_ net185 _04020_ _04021_ net724 vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__a211o_1
X_10787_ _04919_ net505 vssd1 vssd1 vccd1 vccd1 _07127_ sky130_fd_sc_hd__xnor2_1
X_15314_ net1288 vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11260__A1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12526_ net2500 net216 net404 vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__mux2_1
X_16294_ clknet_leaf_92_wb_clk_i _02048_ _00277_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11949__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15245_ net1265 vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12457_ net2380 net190 net411 vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11408_ team_01_WB.instance_to_wrap.cpu.f0.i\[20\] _07700_ _07707_ team_01_WB.instance_to_wrap.cpu.f0.i\[21\]
+ vssd1 vssd1 vccd1 vccd1 _07727_ sky130_fd_sc_hd__a31o_1
X_15176_ net1381 vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__inv_2
X_12388_ net2879 net313 net425 vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08550__C net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14127_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[30\] _04243_ _04254_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[102\]
+ _04412_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__a221o_1
X_11339_ _04469_ _04470_ vssd1 vssd1 vccd1 vccd1 _07668_ sky130_fd_sc_hd__nor2_1
XANTENNA__10771__B1 _07110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09943__A net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14058_ _04217_ _04260_ _04343_ _04346_ _04146_ vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__o41a_1
XANTENNA__11684__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13465__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13009_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[77\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[85\]
+ net864 vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_145_Left_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17817_ clknet_leaf_96_wb_clk_i _03493_ _01757_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[87\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15680__A net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08550_ net1077 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[19\] net901
+ vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__and3_1
X_17748_ clknet_leaf_92_wb_clk_i _03424_ _01688_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16565__CLK clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10320__C net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10826__A1 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08481_ net1029 net885 vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__and2_2
XANTENNA__08495__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17679_ clknet_leaf_127_wb_clk_i _03363_ _01620_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_134_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08294__A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09102_ net1094 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[13\] net910
+ vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_100_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10054__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_154_Left_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09995__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09033_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[9\] net701 _05370_ _05372_
+ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_26_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout308_A _07935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09747__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold310 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1845 sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1856 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold332 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1867 sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1878 sky130_fd_sc_hd__dlygate4sd3_1
Xhold354 _02158_ vssd1 vssd1 vccd1 vccd1 net1889 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12831__X _03650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold365 _01975_ vssd1 vssd1 vccd1 vccd1 net1900 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1911 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10762__B1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold387 net136 vssd1 vssd1 vccd1 vccd1 net1922 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout801 _04646_ vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__buf_6
Xhold398 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1933 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09853__A net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout812 net814 vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__clkbuf_8
X_09935_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[4\] _04634_ net754 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06275_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout823 net824 vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__buf_2
Xfanout834 team_01_WB.instance_to_wrap.cpu.RU0.next_ihit vssd1 vssd1 vccd1 vccd1 net834
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout677_A _04790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout845 net851 vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__clkbuf_2
Xfanout856 net857 vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__clkbuf_4
X_09866_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[12\] net813 net731 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06206_ sky130_fd_sc_hd__a22o_1
Xfanout867 net868 vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10514__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout878 _04810_ vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__clkbuf_8
Xhold1010 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2545 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08469__A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1021 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[16\] vssd1 vssd1 vccd1 vccd1
+ net2556 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout889 net890 vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__buf_4
XANTENNA__09380__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1032 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2567 sky130_fd_sc_hd__dlygate4sd3_1
X_08817_ net1105 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[1\] net942 vssd1
+ vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__and3_1
Xhold1043 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2578 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09291__C net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09797_ net1156 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[14\] net959
+ vssd1 vssd1 vccd1 vccd1 _06137_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_107_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout844_A net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1054 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2589 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout465_X net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1065 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1076 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2611 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15590__A net1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08748_ net1012 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[4\] _04779_
+ vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__and3_1
Xhold1087 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2622 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1098 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2633 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12806__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10230__C net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10817__A1 _05963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_2_0_wb_clk_i_X clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13822__B net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08679_ net1086 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[7\] net904 vssd1
+ vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_124_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ net528 _07049_ _06965_ vssd1 vssd1 vccd1 vccd1 _07050_ sky130_fd_sc_hd__o21ai_1
X_11690_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[13\] _07553_ net717 vssd1 vssd1
+ vccd1 vccd1 _07889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08635__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10641_ _06974_ _06977_ _06978_ net557 vssd1 vssd1 vccd1 vccd1 _06981_ sky130_fd_sc_hd__o22a_1
XANTENNA__11342__B net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10045__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13360_ team_01_WB.instance_to_wrap.cpu.f0.i\[9\] net1070 vssd1 vssd1 vccd1 vccd1
+ _03831_ sky130_fd_sc_hd__xor2_1
XFILLER_0_63_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09986__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10572_ _04746_ _06910_ vssd1 vssd1 vccd1 vccd1 _06912_ sky130_fd_sc_hd__or2_2
X_12311_ net3043 net286 net433 vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__mux2_1
XANTENNA__11769__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13291_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[26\] net825 _03775_ _03777_
+ vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__o22a_1
X_15030_ net1256 vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__inv_2
XANTENNA__14192__B1 net1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12242_ net2316 net229 net441 vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12742__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10979__S1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12173_ net1755 net261 net448 vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11124_ _07451_ _07459_ _07462_ _07463_ vssd1 vssd1 vccd1 vccd1 _07464_ sky130_fd_sc_hd__nor4_1
XFILLER_0_101_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16981_ clknet_leaf_118_wb_clk_i _02668_ _00964_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11055_ net555 _06280_ vssd1 vssd1 vccd1 vccd1 _07395_ sky130_fd_sc_hd__or2_1
X_15932_ net1361 vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__inv_2
XANTENNA__10505__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09371__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10006_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[1\] net809 _06345_ vssd1
+ vssd1 vccd1 vccd1 _06346_ sky130_fd_sc_hd__a21o_1
X_15863_ net1348 vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__inv_2
XANTENNA__09910__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17602_ clknet_leaf_86_wb_clk_i _03289_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_14814_ net1317 vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__inv_2
X_15794_ net1231 vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10808__A1 _07015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17533_ clknet_leaf_66_wb_clk_i _03220_ _01516_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_14745_ net1188 vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__inv_2
X_11957_ net2262 net290 net476 vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17464_ clknet_leaf_38_wb_clk_i _03151_ _01447_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10908_ _06984_ _07000_ net518 vssd1 vssd1 vccd1 vccd1 _07248_ sky130_fd_sc_hd__mux2_1
XANTENNA__10284__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14676_ net1204 vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11888_ net2297 net307 net486 vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09003__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16415_ clknet_leaf_138_wb_clk_i _02169_ _00398_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11252__B _06919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13627_ net186 _04064_ _04065_ net726 vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__a211o_1
X_10839_ _05491_ _06159_ _07177_ _07178_ vssd1 vssd1 vccd1 vccd1 _07179_ sky130_fd_sc_hd__a22oi_2
X_17395_ clknet_leaf_15_wb_clk_i _03082_ _01378_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09426__A1 net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16346_ clknet_leaf_101_wb_clk_i _02100_ _00329_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[69\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__09977__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13558_ net196 net192 _07815_ _07865_ net642 vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__o2111a_1
XPHY_EDGE_ROW_132_Right_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11679__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12509_ net3061 net286 net410 vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__mux2_1
X_16277_ clknet_leaf_125_wb_clk_i _02031_ _00260_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13489_ _03949_ _03843_ vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_89_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18016_ net637 vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_1
X_15228_ net1247 vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12733__A1 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15159_ net1215 vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__inv_2
XANTENNA__10315__C net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09673__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07981_ team_01_WB.instance_to_wrap.cpu.f0.i\[15\] vssd1 vssd1 vccd1 vccd1 _04479_
+ sky130_fd_sc_hd__inv_2
X_09720_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[21\] net820 net818 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__a22o_1
XANTENNA__12303__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09362__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09901__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16279__Q team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09651_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[23\] net786 net776 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08602_ _04920_ _04940_ _04941_ vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__or3_1
X_09582_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[25\] net753 net743 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08533_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[18\] net658 _04853_
+ _04861_ _04864_ vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08295__Y _04635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout258_A _07888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08464_ net1109 net885 vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__and2_2
Xclkbuf_3_7_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_147_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08455__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09417__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08395_ _04708_ _04716_ net712 team_01_WB.instance_to_wrap.cpu.CU0.bit30 vssd1 vssd1
+ vccd1 vccd1 _04735_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout425_A net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1167_A net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09968__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17921__1528 vssd1 vssd1 vccd1 vccd1 net1528 _17921__1528/LO sky130_fd_sc_hd__conb_1
XFILLER_0_115_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout213_X net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08471__B net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1334_A net1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09016_ net1095 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[9\] net930 vssd1
+ vssd1 vccd1 vccd1 _05356_ sky130_fd_sc_hd__and3_1
XANTENNA__14174__B1 net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09286__C net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout794_A net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12724__A1 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold140 net90 vssd1 vssd1 vccd1 vccd1 net1675 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 net100 vssd1 vssd1 vccd1 vccd1 net1686 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 team_01_WB.instance_to_wrap.cpu.f0.write_data\[31\] vssd1 vssd1 vccd1 vccd1
+ net1697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 net1708
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold184 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1719 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 _02012_ vssd1 vssd1 vccd1 vccd1 net1730 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13817__B net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout620 _04846_ vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__buf_2
Xfanout631 _03733_ vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__clkbuf_4
X_09918_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[4\] net796 net736 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06258_ sky130_fd_sc_hd__a22o_1
Xfanout642 net643 vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12213__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout653 _04819_ vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__buf_4
XANTENNA__10522__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout664 _04806_ vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__buf_6
Xfanout675 _04791_ vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09353__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout686 _04778_ vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__buf_8
Xfanout697 net698 vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_126_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09849_ net376 net342 net560 vssd1 vssd1 vccd1 vccd1 _06189_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11160__A0 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout847_X net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12860_ net2111 net292 net380 vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__mux2_1
X_11811_ net2160 net285 net493 vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__mux2_1
XANTENNA__13988__B1 _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09656__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ net1738 net638 net606 _03622_ vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14530_ net1366 vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__inv_2
X_11742_ net1847 net312 net500 vssd1 vssd1 vccd1 vccd1 _03219_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14461_ net1306 vssd1 vssd1 vccd1 vccd1 _00255_ sky130_fd_sc_hd__inv_2
X_11673_ _07812_ _07875_ vssd1 vssd1 vccd1 vccd1 _07876_ sky130_fd_sc_hd__and2b_1
X_16200_ clknet_leaf_158_wb_clk_i _01960_ _00188_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13412_ _04501_ _05224_ vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__or2_1
X_17180_ clknet_leaf_58_wb_clk_i _02867_ _01163_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09959__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10624_ net556 _06858_ _06921_ vssd1 vssd1 vccd1 vccd1 _06964_ sky130_fd_sc_hd__a21o_1
X_14392_ net1186 vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16131_ clknet_leaf_127_wb_clk_i _00022_ _00119_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.state\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13343_ net586 _07688_ _03817_ net828 vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__a31o_1
X_10555_ net545 net513 vssd1 vssd1 vccd1 vccd1 _06895_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14165__B1 net1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16062_ clknet_leaf_154_wb_clk_i _01855_ _00050_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_106_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13274_ net1068 _03754_ vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09196__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10486_ _05870_ _05901_ _05869_ vssd1 vssd1 vccd1 vccd1 _06826_ sky130_fd_sc_hd__o21ba_1
X_15013_ net1286 vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__inv_2
X_12225_ _07794_ _07945_ net573 vssd1 vssd1 vccd1 vccd1 _07962_ sky130_fd_sc_hd__and3_4
XANTENNA__08395__A1 _04708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08395__B2 team_01_WB.instance_to_wrap.cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12156_ net2232 net288 net452 vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__mux2_1
XANTENNA__09924__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11107_ _06905_ _07284_ _07446_ vssd1 vssd1 vccd1 vccd1 _07447_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12123__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16964_ clknet_leaf_83_wb_clk_i _02651_ _00947_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_12087_ net2258 net307 net462 vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_34_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11038_ _07271_ _07272_ vssd1 vssd1 vccd1 vccd1 _07378_ sky130_fd_sc_hd__nand2_1
X_15915_ net1367 vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__inv_2
X_16895_ clknet_leaf_44_wb_clk_i _02582_ _00878_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08698__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11962__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15846_ net1326 vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__inv_2
XANTENNA__08396__X _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13979__B1 _04246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12989_ net2745 net2642 net865 vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__mux2_1
X_15777_ net1197 vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17516_ clknet_leaf_147_wb_clk_i _03203_ _01499_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14728_ net1210 vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14659_ net1306 vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__inv_2
X_17447_ clknet_leaf_99_wb_clk_i _03134_ _01430_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08870__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09668__A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10009__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08180_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[101\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[93\]
+ net1050 vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__mux2_1
X_17378_ clknet_leaf_57_wb_clk_i _03065_ _01361_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13600__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12954__A1 _05074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11710__B net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16329_ clknet_leaf_119_wb_clk_i _02083_ _00312_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[52\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08622__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12822__A net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09583__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10342__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12033__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09690__X _06030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08138__B2 _04483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09335__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09703_ net1154 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[21\] net964
+ vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_71_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11872__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09634_ net1135 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[23\] net968
+ vssd1 vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__and3_1
XANTENNA__08747__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09565_ net1151 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[25\] net969
+ vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__and3_1
XFILLER_0_139_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08466__B net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11445__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08516_ net1077 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[18\] net929
+ vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09496_ _05808_ _05835_ vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08447_ net1109 net919 vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__and2_2
XFILLER_0_147_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout330_X net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout807_A net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout428_X net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11323__D team_01_WB.instance_to_wrap.cpu.DM0.data_i\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11460__X _07756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08482__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08378_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[4\] _04711_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__or3b_1
XFILLER_0_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12208__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08613__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14147__B1 _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10340_ net1139 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[17\] net970
+ vssd1 vssd1 vccd1 vccd1 _06680_ sky130_fd_sc_hd__and3_1
XFILLER_0_143_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout797_X net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12291__X _07964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10271_ net1128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[19\] net948
+ vssd1 vssd1 vccd1 vccd1 _06611_ sky130_fd_sc_hd__and3_1
XFILLER_0_143_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12010_ net3098 net259 net469 vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__mux2_1
XANTENNA__13370__A1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_47_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout964_X net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1404 net1409 vssd1 vssd1 vccd1 vccd1 net1404 sky130_fd_sc_hd__buf_4
Xfanout1415 net1416 vssd1 vssd1 vccd1 vccd1 net1415 sky130_fd_sc_hd__buf_4
Xfanout1426 net1427 vssd1 vssd1 vccd1 vccd1 net1426 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13658__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout450 _07958_ vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09326__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout461 _07955_ vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__clkbuf_8
Xfanout472 _07952_ vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13961_ _04217_ _04220_ _04239_ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__and3_4
XANTENNA__12878__S net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout483 _07948_ vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__clkbuf_8
Xfanout494 _07944_ vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11782__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12912_ net1834 net869 net356 _03683_ vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__a22o_1
X_15700_ net1399 vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__inv_2
X_16680_ clknet_leaf_64_wb_clk_i _02367_ _00663_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09760__B net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12881__A0 team_01_WB.instance_to_wrap.cpu.f0.write_data\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13892_ _04139_ net572 _04197_ vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15631_ net1299 vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_100_Left_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12843_ net1824 net200 net379 vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__mux2_1
XANTENNA__10398__S net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10239__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15562_ net1284 vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__inv_2
X_12774_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] net1061 net362 _03610_
+ vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14513_ net1364 vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__inv_2
X_17301_ clknet_leaf_111_wb_clk_i _02988_ _01284_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11725_ net2256 net277 net502 vssd1 vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_48_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15493_ net1275 vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_859 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14444_ net1224 vssd1 vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__inv_2
X_17232_ clknet_leaf_109_wb_clk_i _02919_ _01215_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11656_ net1992 net242 net501 vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08823__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11739__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13594__D1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10607_ net551 _06280_ vssd1 vssd1 vccd1 vccd1 _06947_ sky130_fd_sc_hd__nor2_1
X_17163_ clknet_leaf_8_wb_clk_i _02850_ _01146_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_86_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14375_ net1208 vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__inv_2
XANTENNA__12118__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11587_ _07803_ vssd1 vssd1 vccd1 vccd1 _07804_ sky130_fd_sc_hd__inv_2
XANTENNA__08604__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16114_ clknet_leaf_136_wb_clk_i _01889_ _00102_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_40_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14138__B1 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13326_ _03798_ _03802_ _03804_ _00020_ vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__a2bb2o_1
Xhold909 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[49\] vssd1 vssd1 vccd1 vccd1
+ net2444 sky130_fd_sc_hd__dlygate4sd3_1
X_17094_ clknet_leaf_72_wb_clk_i _02781_ _01077_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10538_ net1080 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[31\] net906
+ net658 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[31\] vssd1 vssd1 vccd1
+ vccd1 _06878_ sky130_fd_sc_hd__a32o_1
XFILLER_0_12_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12913__Y _03684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11957__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16045_ clknet_leaf_4_wb_clk_i net876 _00033_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.enable
+ sky130_fd_sc_hd__dfrtp_1
X_13257_ net1068 _03748_ vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__or2_1
XANTENNA__13738__A team_01_WB.instance_to_wrap.cpu.DM0.dhit vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10469_ _06798_ _06800_ _06805_ _06808_ vssd1 vssd1 vccd1 vccd1 _06809_ sky130_fd_sc_hd__or4_2
XFILLER_0_86_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12208_ net1858 net258 net445 vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13188_ net21 net835 net628 net1709 vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12139_ net1850 net266 net452 vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10162__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17996_ net635 vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__clkbuf_1
Xhold1609 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net3144 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09951__A net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16947_ clknet_leaf_23_wb_clk_i _02634_ _00930_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13664__A2 _07489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17920__1527 vssd1 vssd1 vccd1 vccd1 net1527 _17920__1527/LO sky130_fd_sc_hd__conb_1
X_16878_ clknet_leaf_38_wb_clk_i _02565_ _00861_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15829_ net1339 vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__inv_2
XANTENNA__11705__B net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08286__B team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09350_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[25\] net678 net653 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[25\]
+ _05686_ vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__a221o_1
X_08301_ net1155 net974 vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__and2_1
X_09281_ net1009 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[22\] net935 vssd1
+ vssd1 vccd1 vccd1 _05621_ sky130_fd_sc_hd__and3_1
XANTENNA__11280__X _07620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08232_ net2381 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[41\] net1057 vssd1 vssd1
+ vccd1 vccd1 _03455_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08163_ net2454 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[110\] net1045 vssd1 vssd1
+ vccd1 vccd1 _03524_ sky130_fd_sc_hd__mux2_1
XANTENNA__12028__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08094_ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[17\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[16\]
+ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[19\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__or4_1
XANTENNA__11867__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload60 clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload60/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload71 clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload71/Y sky130_fd_sc_hd__inv_6
Xclkload82 clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload82/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_141_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1032_A net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload93 clknet_leaf_144_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload93/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_11_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09564__C net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout492_A _07944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10072__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08996_ _05324_ _05327_ net618 net617 vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_110_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12698__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout757_A _04675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11455__X team_01_WB.instance_to_wrap.cpu.DM0.next_enable vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13383__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08477__A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09617_ _05935_ _05954_ _05955_ _05956_ vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__or4_1
XFILLER_0_35_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout924_A _04770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout545_X net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09548_ _05880_ _05885_ _05886_ _05887_ vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__or4_1
XFILLER_0_39_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_120_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14080__A2 _04244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13830__B net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09479_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[30\] net683 _05817_
+ _05818_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__a211o_1
XANTENNA__08924__B net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11510_ net2010 net876 _07758_ _07782_ vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__o22a_1
XFILLER_0_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12490_ net2911 net189 net407 vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__mux2_1
XANTENNA__09739__C net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08643__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12918__A1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11441_ team_01_WB.instance_to_wrap.cpu.f0.i\[6\] _07675_ net324 vssd1 vssd1 vccd1
+ vccd1 _07745_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08047__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14160_ _04195_ _04440_ net1422 vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13591__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11372_ net1072 _07676_ vssd1 vssd1 vccd1 vccd1 _07701_ sky130_fd_sc_hd__nand2_2
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11777__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13111_ net1 net843 vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__nor2_2
XANTENNA__10944__A3 _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10323_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[18\] net745 _06660_ _06661_
+ _06662_ vssd1 vssd1 vccd1 vccd1 _06663_ sky130_fd_sc_hd__a2111o_1
X_14091_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[93\] _04240_ _04263_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[125\]
+ _04377_ vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__a221o_1
XANTENNA__09547__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input53_A wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13042_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[44\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[52\]
+ net858 vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__mux2_1
X_10254_ net339 _06593_ vssd1 vssd1 vccd1 vccd1 _06594_ sky130_fd_sc_hd__nor2_1
XANTENNA__09474__C net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1201 net1207 vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1212 net1223 vssd1 vssd1 vccd1 vccd1 net1212 sky130_fd_sc_hd__clkbuf_4
X_17850_ clknet_leaf_122_wb_clk_i net1758 _01790_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[120\]
+ sky130_fd_sc_hd__dfrtp_1
X_10185_ _06517_ _06521_ _06523_ _06524_ vssd1 vssd1 vccd1 vccd1 _06525_ sky130_fd_sc_hd__a31o_2
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1223 net1304 vssd1 vssd1 vccd1 vccd1 net1223 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08770__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10413__C net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1234 net1235 vssd1 vssd1 vccd1 vccd1 net1234 sky130_fd_sc_hd__buf_2
X_16801_ clknet_leaf_56_wb_clk_i _02488_ _00784_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1245 net1248 vssd1 vssd1 vccd1 vccd1 net1245 sky130_fd_sc_hd__clkbuf_4
Xfanout1256 net1258 vssd1 vssd1 vccd1 vccd1 net1256 sky130_fd_sc_hd__buf_4
Xfanout1267 net1268 vssd1 vssd1 vccd1 vccd1 net1267 sky130_fd_sc_hd__buf_2
X_17781_ clknet_leaf_95_wb_clk_i _03457_ _01721_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[51\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout280 net283 vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__buf_2
X_14993_ net1419 vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__inv_2
Xfanout1278 net1281 vssd1 vssd1 vccd1 vccd1 net1278 sky130_fd_sc_hd__buf_4
Xfanout291 _07941_ vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__clkbuf_2
Xfanout1289 net1302 vssd1 vssd1 vccd1 vccd1 net1289 sky130_fd_sc_hd__buf_2
X_16732_ clknet_leaf_60_wb_clk_i _02419_ _00715_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12401__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13944_ _04225_ _04234_ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__nor2_4
XANTENNA__08818__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13875_ _04184_ _04185_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[11\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__a211o_1
X_16663_ clknet_leaf_14_wb_clk_i _02350_ _00646_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12826_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[2\] _07489_ net1037 vssd1 vssd1
+ vccd1 vccd1 _03647_ sky130_fd_sc_hd__mux2_1
X_15614_ net1317 vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__inv_2
X_16594_ clknet_leaf_143_wb_clk_i _02281_ _00577_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14071__A2 _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12757_ net1585 net638 net607 _03599_ vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__a22o_1
X_15545_ net1236 vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10093__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11708_ net612 _07804_ _07903_ _07902_ vssd1 vssd1 vccd1 vccd1 _07904_ sky130_fd_sc_hd__a31o_4
XFILLER_0_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15476_ net1378 vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__inv_2
X_12688_ net3036 net189 net383 vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__mux2_1
XANTENNA__09011__A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17215_ clknet_leaf_41_wb_clk_i _02902_ _01198_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14427_ net1325 vssd1 vssd1 vccd1 vccd1 _00221_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11639_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[24\] net713 net616 vssd1 vssd1
+ vccd1 vccd1 _07849_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10157__A net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13582__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17146_ clknet_leaf_76_wb_clk_i _02833_ _01129_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09946__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14358_ net1333 vssd1 vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold706 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 net2241
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold717 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold728 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2263 sky130_fd_sc_hd__dlygate4sd3_1
X_13309_ _07686_ _07709_ _03790_ net587 vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_94_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17077_ clknet_leaf_110_wb_clk_i _02764_ _01060_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold739 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2274 sky130_fd_sc_hd__dlygate4sd3_1
X_14289_ net1346 vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13334__A1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16028_ net1335 vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_90_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08850_ net599 _05187_ _05188_ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__o21a_2
XANTENNA__15683__A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1406 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2941 sky130_fd_sc_hd__dlygate4sd3_1
X_08781_ net1094 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[0\] net922 vssd1
+ vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__and3_1
Xhold1417 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[90\] vssd1 vssd1 vccd1 vccd1
+ net2952 sky130_fd_sc_hd__dlygate4sd3_1
X_17979_ net1494 vssd1 vssd1 vccd1 vccd1 la_data_out[21] sky130_fd_sc_hd__buf_2
Xhold1428 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2963 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17671__Q team_01_WB.instance_to_wrap.cpu.DM0.readdata\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1439 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[19\] vssd1 vssd1 vccd1 vccd1
+ net2974 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11648__A1 _07154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11716__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12311__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_140_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09402_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[27\] net672 net667 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[27\]
+ _05738_ vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_49_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09069__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10871__A2 _06032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14062__A2 _04245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08277__A0 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09333_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[24\] net663 net659 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_3_7_0_wb_clk_i_X clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10766__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout240_A _07870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout338_A _06903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10084__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09264_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[20\] net665 net652 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[20\]
+ _05603_ vssd1 vssd1 vccd1 vccd1 _05604_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08215_ net2432 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[58\] net1052 vssd1 vssd1
+ vccd1 vccd1 _03472_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09195_ net1004 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[17\] net923 vssd1
+ vssd1 vccd1 vccd1 _05535_ sky130_fd_sc_hd__and3_1
XANTENNA__10067__A _06280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout505_A _06636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1247_A net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09777__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08146_ _04580_ _04581_ _04586_ _04587_ _04584_ vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__o221a_1
XFILLER_0_114_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09241__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08077_ _04515_ _04538_ _04544_ vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_112_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1035_X net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1414_A net1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13097__B net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09294__C net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout874_A net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout495_X net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold11 _02015_ vssd1 vssd1 vccd1 vccd1 net1546 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[18\] vssd1 vssd1 vccd1 vccd1 net1557
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 net146 vssd1 vssd1 vccd1 vccd1 net1568 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13825__B net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08979_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[8\] net688 _05316_ _05317_
+ _05318_ vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__a2111oi_1
Xhold44 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[16\] vssd1 vssd1 vccd1 vccd1 net1579
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout662_X net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold55 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[26\] vssd1 vssd1 vccd1 vccd1
+ net1590 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13628__A2 _07269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08919__B _05224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold66 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1 net1601
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 _01985_ vssd1 vssd1 vccd1 vccd1 net1612 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12221__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold88 _02005_ vssd1 vssd1 vccd1 vccd1 net1623 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ net1927 net315 net473 vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__mux2_1
Xhold99 team_01_WB.instance_to_wrap.a1.ADR_I\[11\] vssd1 vssd1 vccd1 vccd1 net1634
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08504__A1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08638__C net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11103__A3 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10941_ net527 _07280_ _07150_ _07062_ vssd1 vssd1 vccd1 vccd1 _07281_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_98_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout927_X net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13660_ net989 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] _04091_ _04092_
+ vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10872_ _07210_ _07211_ net519 vssd1 vssd1 vccd1 vccd1 _07212_ sky130_fd_sc_hd__mux2_1
X_12611_ net2695 net282 net398 vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13591_ net721 _07611_ net1074 vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_27_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10676__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11361__A team_01_WB.instance_to_wrap.cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_54_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15330_ net1320 vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__inv_2
X_12542_ net1880 net284 net405 vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09469__C net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09480__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15261_ net1236 vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12473_ net2510 net229 net413 vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__mux2_1
X_17000_ clknet_leaf_64_wb_clk_i _02687_ _00983_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_14212_ net1566 vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13564__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11424_ _04485_ _07701_ vssd1 vssd1 vccd1 vccd1 _07736_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09768__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15192_ net1212 vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09232__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_8 _03654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14143_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[103\] _04254_ _04264_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[111\]
+ _04427_ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__a221o_1
X_11355_ _04484_ _07683_ vssd1 vssd1 vccd1 vccd1 _07684_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10306_ _06642_ _06643_ _06644_ _06645_ vssd1 vssd1 vccd1 vccd1 _06646_ sky130_fd_sc_hd__or4_1
X_14074_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[36\] _04230_ _04251_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[84\]
+ _04361_ vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__a221o_1
X_11286_ _07019_ _07056_ _07111_ vssd1 vssd1 vccd1 vccd1 _07626_ sky130_fd_sc_hd__or3_1
X_17902_ net1437 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
X_13025_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[61\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[69\]
+ net859 vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__mux2_1
X_10237_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[9\] net803 net749 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06577_ sky130_fd_sc_hd__a22o_1
XANTENNA__11878__A1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1020 net1021 vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__clkbuf_2
Xfanout1031 _04490_ vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__buf_2
XANTENNA__09940__B1 _06278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1042 net1059 vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__clkbuf_4
X_17833_ clknet_leaf_96_wb_clk_i _03509_ _01773_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[103\]
+ sky130_fd_sc_hd__dfrtp_1
X_10168_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[10\] net820 _06506_
+ _06507_ vssd1 vssd1 vccd1 vccd1 _06508_ sky130_fd_sc_hd__a211o_1
Xfanout1053 net1058 vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__clkbuf_2
Xfanout1064 net1065 vssd1 vssd1 vccd1 vccd1 net1064 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_156_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1075 net1076 vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__clkbuf_2
Xfanout1086 net1088 vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15008__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17764_ clknet_leaf_91_wb_clk_i net2213 _01704_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12827__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12131__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1097 net1103 vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__buf_2
XFILLER_0_89_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10099_ _05264_ _05265_ _05301_ net377 vssd1 vssd1 vccd1 vccd1 _06439_ sky130_fd_sc_hd__o31a_1
X_14976_ net1238 vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_63_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08548__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16715_ clknet_leaf_9_wb_clk_i _02402_ _00698_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13927_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[2\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__and2b_2
XFILLER_0_156_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17695_ clknet_leaf_137_wb_clk_i _03379_ _01636_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13868__A_N net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11970__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16646_ clknet_leaf_90_wb_clk_i _02333_ _00629_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13858_ net1180 net1067 net2132 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[19\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14044__A2 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12809_ net364 _03633_ _03634_ net1062 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__a32o_1
X_16577_ clknet_leaf_57_wb_clk_i _02264_ _00560_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10439__X _06779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13252__B1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13789_ _04154_ _04171_ _04172_ _04167_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__a31o_1
XFILLER_0_32_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15528_ net1382 vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_44_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12654__X _03569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15459_ net1270 vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08000_ team_01_WB.instance_to_wrap.cpu.f0.num\[2\] vssd1 vssd1 vccd1 vccd1 _04498_
+ sky130_fd_sc_hd__inv_2
XANTENNA__13555__A1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12814__B _07507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold503 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2038 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16570__Q team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17129_ clknet_leaf_36_wb_clk_i _02816_ _01112_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold514 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2049 sky130_fd_sc_hd__dlygate4sd3_1
Xhold525 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2060 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12306__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold536 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2071 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13307__A1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold547 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[3\] vssd1 vssd1 vccd1 vccd1
+ net2082 sky130_fd_sc_hd__dlygate4sd3_1
X_09951_ net1155 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[3\] net959 vssd1
+ vssd1 vccd1 vccd1 _06291_ sky130_fd_sc_hd__and3_1
Xhold558 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2093 sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2104 sky130_fd_sc_hd__dlygate4sd3_1
X_08902_ net1108 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[2\] net898 vssd1
+ vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__and3_1
XFILLER_0_148_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09882_ net1152 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[5\] net957 vssd1
+ vssd1 vccd1 vccd1 _06222_ sky130_fd_sc_hd__and3_1
XANTENNA__08579__X _04919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09931__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08833_ net1105 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[1\] net915 vssd1
+ vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__and3_1
XANTENNA__08734__B2 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[5\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1203 _03460_ vssd1 vssd1 vccd1 vccd1 net2738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1214 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2749 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1225 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2760 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout288_A _07941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1236 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[87\] vssd1 vssd1 vccd1 vccd1
+ net2771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1247 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2782 sky130_fd_sc_hd__dlygate4sd3_1
X_08764_ _05100_ _05101_ _05102_ _05103_ vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__or4_1
XANTENNA__12041__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1258 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[114\] vssd1 vssd1 vccd1 vccd1
+ net2793 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1269 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2804 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08458__C net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12294__A1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08695_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[7\] net656 _05014_ _05021_
+ _05024_ vssd1 vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout455_A _07956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11880__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1197_A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_146_Right_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08755__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout622_A net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09316_ net1121 net711 net600 net594 vssd1 vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11254__C1 _06903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09998__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09289__C net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09247_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[21\] net700 _05586_ net706
+ vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout410_X net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1152_X net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout508_X net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09178_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[16\] net690 _05515_ _05516_
+ _05517_ vssd1 vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_16_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09214__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08129_ _04470_ team_01_WB.instance_to_wrap.cpu.f0.num\[25\] team_01_WB.instance_to_wrap.cpu.f0.num\[15\]
+ _04479_ _04598_ vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12216__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11140_ net334 net337 _07390_ vssd1 vssd1 vccd1 vccd1 _07480_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout877_X net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__buf_2
X_11071_ _07409_ _07410_ _07373_ vssd1 vssd1 vccd1 vccd1 _07411_ sky130_fd_sc_hd__a21bo_1
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__buf_2
X_10022_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[1\] net740 _06359_ _06360_
+ _06361_ vssd1 vssd1 vccd1 vccd1 _06362_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11356__A _04483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14830_ net1299 vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_129_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12809__B1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input16_A DAT_I[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14761_ net1283 vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__inv_2
X_11973_ net2242 net236 net471 vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__mux2_1
XANTENNA__13482__B1 _05705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11790__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12824__A3 _03645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16500_ clknet_leaf_156_wb_clk_i _02254_ _00483_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10296__B1 _06634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13712_ net1548 _04504_ _03573_ vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__a21bo_1
X_10924_ net328 _07263_ _07262_ _07260_ vssd1 vssd1 vccd1 vccd1 _07264_ sky130_fd_sc_hd__a211o_1
X_17480_ clknet_leaf_27_wb_clk_i _03167_ _01463_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_14692_ net1195 vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14026__A2 _04244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16431_ clknet_leaf_139_wb_clk_i _02185_ _00414_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10855_ net376 net330 vssd1 vssd1 vccd1 vccd1 _07195_ sky130_fd_sc_hd__nor2_1
X_13643_ net187 _04077_ _04078_ net725 vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__a211o_1
XFILLER_0_67_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08384__B net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10048__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16362_ clknet_leaf_101_wb_clk_i _02116_ _00345_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[85\]
+ sky130_fd_sc_hd__dfstp_1
X_13574_ net196 net192 _07876_ net642 vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__o211a_1
XANTENNA__09199__C net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10786_ _04919_ net505 net369 vssd1 vssd1 vccd1 vccd1 _07126_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09453__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15313_ net1393 vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__inv_2
XANTENNA__08378__C_N team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12525_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[29\] net220 net404 vssd1
+ vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16293_ clknet_leaf_123_wb_clk_i _02047_ _00276_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15244_ net1257 vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__inv_2
X_12456_ _07790_ _07946_ net573 vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_10_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_110_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_110_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_140_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08831__C net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11407_ _07712_ _07726_ vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__nor2_1
X_15175_ net1390 vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__inv_2
X_12387_ net2095 net317 net426 vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12126__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14126_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[78\] _04235_ _04241_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[94\]
+ vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11338_ _07667_ net1985 _07655_ vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__mux2_1
XANTENNA__10771__A1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11965__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14057_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\] _04237_ _04342_ _04344_
+ _04345_ vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__a2111o_1
X_11269_ net338 _06959_ vssd1 vssd1 vccd1 vccd1 _07609_ sky130_fd_sc_hd__nand2_1
X_13008_ net2912 net2878 net854 vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__mux2_1
X_17816_ clknet_leaf_120_wb_clk_i net2747 _01756_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[86\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_89_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17747_ clknet_leaf_92_wb_clk_i _03423_ _01687_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14959_ net1386 vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__inv_2
XANTENNA__10287__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08480_ net1081 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[23\] net897
+ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__and3_1
X_17678_ clknet_leaf_157_wb_clk_i net1171 _01619_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.pc_enable
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14017__A2 _04236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09692__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16629_ clknet_leaf_112_wb_clk_i _02316_ _00612_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08294__B net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11236__C1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09101_ net1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[13\] net914
+ vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__and3_1
XFILLER_0_57_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09032_ _05363_ _05364_ _05365_ _05371_ vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__or4_2
XANTENNA__13528__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11539__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08741__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold300 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[28\] vssd1 vssd1 vccd1 vccd1 net1835
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[27\] vssd1 vssd1 vccd1 vccd1 net1846
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12036__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10345__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout203_A _07855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold322 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1857 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10211__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold333 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1868 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold344 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1890 sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1901 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11875__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold377 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1912 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout802 _04643_ vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__clkbuf_8
Xhold388 _01972_ vssd1 vssd1 vccd1 vccd1 net1923 sky130_fd_sc_hd__dlygate4sd3_1
X_09934_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[4\] net815 net738 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06274_ sky130_fd_sc_hd__a22o_1
Xhold399 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1934 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout813 net814 vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1112_A net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout824 _04630_ vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__clkbuf_4
Xfanout835 _03737_ vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__clkbuf_4
Xfanout846 net847 vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__buf_2
X_09865_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[12\] net792 net789 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06205_ sky130_fd_sc_hd__a22o_1
XANTENNA_input8_A DAT_I[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout857 net858 vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__clkbuf_4
Xhold1000 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2535 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09572__C net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11711__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout868 _03718_ vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__clkbuf_2
Xhold1011 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2546 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout879 _04810_ vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__buf_2
Xhold1022 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2557 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1033 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[87\] vssd1 vssd1 vccd1 vccd1
+ net2568 sky130_fd_sc_hd__dlygate4sd3_1
X_08816_ net1104 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[1\] net920 vssd1
+ vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__and3_1
X_09796_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[14\] net819 net751 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06136_ sky130_fd_sc_hd__a22o_1
Xhold1044 team_01_WB.instance_to_wrap.cpu.f0.num\[3\] vssd1 vssd1 vccd1 vccd1 net2579
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1055 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2590 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1066 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2601 sky130_fd_sc_hd__dlygate4sd3_1
X_08747_ net1099 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[4\] net893 vssd1
+ vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__and3_1
Xhold1077 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2612 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17635__CLK clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout360_X net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1088 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1099 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2634 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout458_X net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout837_A _03736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13391__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08678_ net1006 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[7\] net911 vssd1
+ vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_124_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10817__A2 _06779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14008__A2 _04258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09683__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout625_X net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10640_ net522 _06928_ vssd1 vssd1 vccd1 vccd1 _06980_ sky130_fd_sc_hd__nand2_1
XANTENNA__08772__X _05112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09435__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_971 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11242__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10571_ _04746_ _06910_ vssd1 vssd1 vccd1 vccd1 _06911_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12310_ net2968 net255 net432 vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__mux2_1
XANTENNA__13519__A1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13290_ net566 _03752_ _03776_ net828 vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout994_X net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08651__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12727__C1 net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12241_ net1977 net261 net440 vssd1 vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__mux2_1
XANTENNA__10255__A net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12742__A2 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12172_ net2320 net267 net447 vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11785__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11123_ _05261_ _06957_ _07101_ vssd1 vssd1 vccd1 vccd1 _07463_ sky130_fd_sc_hd__and3_1
XFILLER_0_130_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10542__X _06882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16980_ clknet_leaf_21_wb_clk_i _02667_ _00963_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11054_ _07062_ _07385_ _07391_ _07392_ _07393_ vssd1 vssd1 vccd1 vccd1 _07394_ sky130_fd_sc_hd__a311o_1
X_15931_ net1367 vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__inv_2
XANTENNA__08379__B team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10005_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[1\] net783 net743 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06345_ sky130_fd_sc_hd__a22o_1
X_15862_ net1345 vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__inv_2
XANTENNA__10421__C net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17601_ clknet_leaf_86_wb_clk_i _03288_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_14813_ net1311 vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__inv_2
X_15793_ net1231 vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__inv_2
X_17532_ clknet_leaf_58_wb_clk_i _03219_ _01515_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14744_ net1191 vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__inv_2
X_11956_ net2012 net316 net477 vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08826__C net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10907_ net375 _06934_ _07014_ _07246_ vssd1 vssd1 vccd1 vccd1 _07247_ sky130_fd_sc_hd__a31o_1
XANTENNA__13207__B1 _03738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17463_ clknet_leaf_13_wb_clk_i _03150_ _01446_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11887_ net2546 net311 net486 vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__mux2_1
X_14675_ net1225 vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_15_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16414_ clknet_leaf_124_wb_clk_i _02168_ _00397_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10838_ _05491_ net330 _07176_ net335 _06915_ vssd1 vssd1 vccd1 vccd1 _07178_ sky130_fd_sc_hd__o221a_1
X_13626_ net199 net195 _07802_ _07907_ net645 vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__o2111a_1
X_17394_ clknet_leaf_110_wb_clk_i _03081_ _01377_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16345_ clknet_leaf_118_wb_clk_i _02099_ _00328_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[68\]
+ sky130_fd_sc_hd__dfstp_1
X_13557_ _03925_ _04006_ vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10769_ net556 _07107_ _07108_ _06963_ vssd1 vssd1 vccd1 vccd1 _07109_ sky130_fd_sc_hd__o22a_1
XFILLER_0_82_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12508_ net2096 net253 net408 vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__mux2_1
X_16276_ clknet_leaf_88_wb_clk_i _00004_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[5\]
+ sky130_fd_sc_hd__dfxtp_4
X_13488_ _03844_ _03845_ _03946_ _05780_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__a32o_1
X_18015_ net637 vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08561__C net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15227_ net1255 vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__inv_2
X_12439_ net2369 net261 net416 vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09954__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15158_ net1256 vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_39_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14109_ _04348_ _04395_ _04376_ net1183 vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__o211a_1
X_15089_ net1423 vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__inv_2
X_07980_ team_01_WB.instance_to_wrap.cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1 _04478_
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_56_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09650_ _05986_ _05987_ _05988_ _05989_ vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__or4_1
X_08601_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[15\] net694 net650 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__a22o_1
X_09581_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[25\] net795 _05905_ _05907_
+ _05912_ vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_89_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09114__A1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08532_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[18\] net699 _04854_ _04860_
+ _04862_ vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_148_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08463_ net1116 net1119 net1125 net1122 vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__nor4b_2
XFILLER_0_77_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08394_ net1170 _04717_ vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__nand2_1
XANTENNA__10059__B _06398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout320_A _07937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08625__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout418_A _03562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1062_A team_01_WB.instance_to_wrap.cpu.RU0.state\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire962_X net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10432__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09567__C net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09015_ net1013 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[9\] net905 vssd1
+ vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__and3_1
XANTENNA__10075__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1327_A net1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold130 team_01_WB.instance_to_wrap.cpu.f0.write_data\[17\] vssd1 vssd1 vccd1 vccd1
+ net1665 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_37_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold141 _02021_ vssd1 vssd1 vccd1 vccd1 net1676 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold152 _02001_ vssd1 vssd1 vccd1 vccd1 net1687 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 _01832_ vssd1 vssd1 vccd1 vccd1 net1698 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10735__B2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold174 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 net1709
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold185 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[9\] vssd1 vssd1 vccd1 vccd1
+ net1720 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10803__A _05657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold196 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[27\] vssd1 vssd1 vccd1 vccd1
+ net1731 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout610 _07685_ vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1115_X net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09917_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[4\] net787 net776 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[4\]
+ _06256_ vssd1 vssd1 vccd1 vccd1 _06257_ sky130_fd_sc_hd__a221o_1
Xfanout632 _03733_ vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__clkbuf_2
Xfanout643 _04839_ vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout954_A net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout654 _04817_ vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout665 _04804_ vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__buf_6
Xfanout676 _04790_ vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_13_Left_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout687 _04776_ vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__buf_6
X_09848_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] net625 _06186_ _06187_
+ vssd1 vssd1 vccd1 vccd1 _06188_ sky130_fd_sc_hd__a22o_2
Xfanout698 _04763_ vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_126_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11160__A1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout742_X net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13833__B net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09779_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[15\] net795 net743 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11810_ net2665 net254 net492 vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] net1060 net362 _03621_
+ vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09656__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08646__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11741_ _07927_ _07928_ _07930_ net613 vssd1 vssd1 vccd1 vccd1 _07931_ sky130_fd_sc_hd__a22o_2
XANTENNA__11463__A2 _07755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11672_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\]
+ _07809_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] vssd1 vssd1 vccd1 vccd1
+ _07875_ sky130_fd_sc_hd__a31o_1
X_14460_ net1228 vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__inv_2
XANTENNA__09408__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10623_ net557 _06858_ _06921_ vssd1 vssd1 vccd1 vccd1 _06963_ sky130_fd_sc_hd__a21oi_4
X_13411_ _03870_ _03871_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__and2b_1
XFILLER_0_153_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14391_ net1186 vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__inv_2
XANTENNA__08616__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_76_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_12__f_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13342_ _04481_ _07687_ vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__nand2_1
X_16130_ clknet_leaf_126_wb_clk_i _00021_ _00118_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10423__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10554_ _06890_ _06893_ net519 vssd1 vssd1 vccd1 vccd1 _06894_ sky130_fd_sc_hd__mux2_1
XANTENNA__12963__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10974__B2 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16061_ clknet_leaf_154_wb_clk_i _01854_ _00049_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\]
+ sky130_fd_sc_hd__dfrtp_4
X_13273_ _03749_ _03762_ vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10485_ _06750_ _06819_ _06823_ _05902_ vssd1 vssd1 vccd1 vccd1 _06825_ sky130_fd_sc_hd__a211o_1
XFILLER_0_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12224_ _07784_ _07789_ _07960_ vssd1 vssd1 vccd1 vccd1 _07961_ sky130_fd_sc_hd__and3_1
X_15012_ net1220 vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__inv_2
XANTENNA__10416__C net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10726__A1 _05898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12155_ net2966 net314 net453 vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__mux2_1
XANTENNA__12404__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11106_ net375 _07330_ _07445_ net531 vssd1 vssd1 vccd1 vccd1 _07446_ sky130_fd_sc_hd__a22o_1
X_12086_ net1951 net309 net460 vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__mux2_1
X_16963_ clknet_leaf_23_wb_clk_i _02650_ _00946_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13676__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11037_ _07375_ _07376_ _07374_ vssd1 vssd1 vccd1 vccd1 _07377_ sky130_fd_sc_hd__a21oi_1
X_15914_ net1352 vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__inv_2
X_16894_ clknet_leaf_85_wb_clk_i _02581_ _00877_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09895__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15845_ net1325 vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15776_ net1197 vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12988_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[98\] net2772 net864 vssd1 vssd1
+ vccd1 vccd1 _02137_ sky130_fd_sc_hd__mux2_1
XANTENNA__09647__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09014__A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17515_ clknet_leaf_7_wb_clk_i _03202_ _01498_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08556__C net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14727_ net1210 vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11939_ net1807 net234 net475 vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10662__A0 _06526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17446_ clknet_leaf_83_wb_clk_i _03133_ _01429_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09949__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14658_ net1224 vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08607__A0 _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13609_ net989 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] _04049_ _04050_
+ vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__a22o_1
X_17377_ clknet_leaf_56_wb_clk_i _03064_ _01360_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14589_ net1412 vssd1 vssd1 vccd1 vccd1 _00383_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16328_ clknet_leaf_95_wb_clk_i _02082_ _00311_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10965__A1 _05263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10607__B _06280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15686__A net1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16259_ clknet_leaf_152_wb_clk_i net1605 _00247_ vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10326__C net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17674__Q team_01_WB.instance_to_wrap.cpu.DM0.readdata\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12314__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09971__X _06311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13131__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09702_ net1145 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[21\] net978
+ vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_71_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10910__X _07250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11142__A1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09633_ net993 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[23\] net951 vssd1
+ vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__and3_1
XANTENNA__12890__A1 _03667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout270_A _07866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09564_ net1149 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[25\] net985
+ vssd1 vssd1 vccd1 vccd1 _05904_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_4_8__f_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14092__B1 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08515_ net1078 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[18\] net878
+ vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_110_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_148_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09495_ _05833_ _05834_ net597 vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__mux2_4
XFILLER_0_78_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout535_A _05190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1277_A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11741__X _07931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08446_ net1083 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[23\] net906
+ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__and3_1
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13198__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08377_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[4\] _04711_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__nor3b_2
XANTENNA_fanout702_A _04758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1065_X net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12945__A2 _03705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09271__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09297__C net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09810__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15596__A net1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09594__A net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10270_ net1128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[19\] net981
+ vssd1 vssd1 vccd1 vccd1 _06610_ sky130_fd_sc_hd__and3_1
XFILLER_0_143_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13828__B net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10708__A1 _06912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout692_X net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1405 net1409 vssd1 vssd1 vccd1 vccd1 net1405 sky130_fd_sc_hd__clkbuf_4
Xfanout1416 net1428 vssd1 vssd1 vccd1 vccd1 net1416 sky130_fd_sc_hd__buf_2
Xfanout1427 net1428 vssd1 vssd1 vccd1 vccd1 net1427 sky130_fd_sc_hd__clkbuf_4
Xfanout440 _07962_ vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08003__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout957_X net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13122__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout451 _07957_ vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__clkbuf_8
Xfanout462 _07955_ vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__buf_4
X_13960_ _04217_ _04220_ _04223_ vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_6_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout473 _07952_ vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__buf_6
Xfanout484 _07948_ vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08497__X _04837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11133__B2 _06919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout495 net498 vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__buf_6
X_12911_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[19\] _03682_ net1036 vssd1
+ vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__mux2_1
X_13891_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[0\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__or2_1
X_15630_ net1297 vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__inv_2
XANTENNA__10892__B1 _07230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12842_ net2749 net205 net379 vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__mux2_1
XANTENNA__14083__B1 _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15561_ net1295 vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__inv_2
X_12773_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[18\] _07251_ net1033 vssd1 vssd1
+ vccd1 vccd1 _03610_ sky130_fd_sc_hd__mux2_1
XANTENNA__08837__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17353__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17300_ clknet_leaf_21_wb_clk_i _02987_ _01283_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14512_ net1353 vssd1 vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11724_ _07913_ _07914_ _07916_ net614 vssd1 vssd1 vccd1 vccd1 _07917_ sky130_fd_sc_hd__a22o_2
XFILLER_0_127_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15492_ net1233 vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13189__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11370__Y _07699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17231_ clknet_leaf_34_wb_clk_i _02918_ _01214_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11655_ net611 _07816_ _07861_ _07860_ vssd1 vssd1 vccd1 vccd1 _07862_ sky130_fd_sc_hd__a31o_2
X_14443_ net1224 vssd1 vssd1 vccd1 vccd1 _00237_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_88_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10606_ net547 _06250_ vssd1 vssd1 vccd1 vccd1 _06946_ sky130_fd_sc_hd__nor2_1
X_17162_ clknet_leaf_32_wb_clk_i _02849_ _01145_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08960__X _05300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11586_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\]
+ _07801_ vssd1 vssd1 vccd1 vccd1 _07803_ sky130_fd_sc_hd__and3_1
X_14374_ net1208 vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09801__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16113_ clknet_leaf_136_wb_clk_i _01888_ _00101_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[20\]
+ sky130_fd_sc_hd__dfrtp_4
X_13325_ _07705_ _03803_ net826 vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__o21ai_1
X_10537_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[31\] net662 net652 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[31\]
+ _06876_ vssd1 vssd1 vccd1 vccd1 _06877_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_17_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09000__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17093_ clknet_leaf_47_wb_clk_i _02780_ _01076_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16044_ clknet_leaf_88_wb_clk_i _01838_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13256_ team_01_WB.instance_to_wrap.cpu.f0.i\[26\] _03747_ vssd1 vssd1 vccd1 vccd1
+ _03748_ sky130_fd_sc_hd__or2_1
X_10468_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[26\] net795 net770 _06806_
+ _06807_ vssd1 vssd1 vccd1 vccd1 _06808_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12207_ net2439 net229 net445 vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__mux2_1
XANTENNA__12134__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13187_ net22 net835 net628 net1668 vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__o22a_1
X_10399_ _05529_ _05730_ vssd1 vssd1 vccd1 vccd1 _06739_ sky130_fd_sc_hd__xor2_1
XANTENNA__10175__A2 _04659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17997__1506 vssd1 vssd1 vccd1 vccd1 _17997__1506/HI net1506 sky130_fd_sc_hd__conb_1
XANTENNA__09009__A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12138_ net2048 net233 net451 vssd1 vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__mux2_1
X_17995_ net637 vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__clkbuf_1
XANTENNA__13649__B1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10162__B net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09317__A1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11973__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13113__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11826__X _07947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08997__A1_N team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[8\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16946_ clknet_leaf_110_wb_clk_i _02633_ _00929_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_12069_ net3132 net241 net461 vssd1 vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__mux2_1
XANTENNA__08848__A net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09670__C net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12872__A1 _03654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16877_ clknet_leaf_67_wb_clk_i _02564_ _00860_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15828_ net1339 vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__inv_2
XANTENNA__14074__B1 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15759_ net1342 vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__inv_2
X_08300_ net1166 net1165 net1161 net1159 vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__and4b_4
XFILLER_0_74_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09280_ _05595_ _05619_ vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08583__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08231_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[50\] net2372 net1053 vssd1 vssd1
+ vccd1 vccd1 _03456_ sky130_fd_sc_hd__mux2_1
XANTENNA__16573__Q team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17429_ clknet_leaf_112_wb_clk_i _03116_ _01412_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12309__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08162_ net2709 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[111\] net1048 vssd1 vssd1
+ vccd1 vccd1 _03525_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08093_ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[21\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[20\]
+ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[23\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload50 clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload50/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA_clkbuf_4_11__f_wb_clk_i_X clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkload61 clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload61/Y sky130_fd_sc_hd__bufinv_16
Xclkload72 clknet_leaf_55_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload72/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload83 clknet_leaf_139_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload83/Y sky130_fd_sc_hd__inv_6
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload94 clknet_leaf_145_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload94/Y sky130_fd_sc_hd__inv_6
XANTENNA__08359__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12044__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1025_A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10166__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_145_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08995_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[8\] net664 _05332_ _05333_
+ _05334_ vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__11883__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout485_A _07948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08758__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09859__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11115__B2 _05263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13383__B _05780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout652_A _04819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1394_A net1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08477__B net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10874__A0 _05898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08531__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09616_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[24\] net740 _05937_ _05943_
+ _05948_ vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout440_X net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09547_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[28\] net785 net761 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout917_A net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09478_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[30\] net664 net650 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08924__C net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08429_ net1081 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[23\] net925
+ vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__and3_1
XANTENNA__12219__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout705_X net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11440_ net324 _07701_ _07744_ vssd1 vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__and3_1
XANTENNA__09876__X _06216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload0 clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload0/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_135_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08047__B2 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10929__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08598__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11371_ net1071 team_01_WB.instance_to_wrap.cpu.f0.i\[6\] _07675_ vssd1 vssd1 vccd1
+ vccd1 _07700_ sky130_fd_sc_hd__and3_2
XFILLER_0_34_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13328__C1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13110_ team_01_WB.instance_to_wrap.a1.curr_state\[2\] team_01_WB.instance_to_wrap.a1.curr_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__or2_1
X_10322_ net1129 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[18\] net975
+ vssd1 vssd1 vccd1 vccd1 _06662_ sky130_fd_sc_hd__and3_1
X_14090_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[45\] _04256_ _04264_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[109\]
+ vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13041_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[45\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[53\]
+ net859 vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__mux2_1
X_10253_ _05374_ _06592_ vssd1 vssd1 vccd1 vccd1 _06593_ sky130_fd_sc_hd__xnor2_2
X_10184_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[10\] net766 vssd1 vssd1
+ vccd1 vccd1 _06524_ sky130_fd_sc_hd__nor2_1
Xfanout1202 net1203 vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__buf_4
XANTENNA_input46_A wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1213 net1216 vssd1 vssd1 vccd1 vccd1 net1213 sky130_fd_sc_hd__buf_4
Xfanout1224 net1226 vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__buf_4
XANTENNA__11793__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16800_ clknet_leaf_45_wb_clk_i _02487_ _00783_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11646__X _07855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1235 net1242 vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__buf_4
XANTENNA__08770__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1246 net1247 vssd1 vssd1 vccd1 vccd1 net1246 sky130_fd_sc_hd__buf_4
X_17780_ clknet_leaf_91_wb_clk_i net2373 _01720_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[50\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1257 net1258 vssd1 vssd1 vccd1 vccd1 net1257 sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_135_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_135_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11106__A1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14992_ net1272 vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__inv_2
Xfanout1268 net1269 vssd1 vssd1 vccd1 vccd1 net1268 sky130_fd_sc_hd__buf_2
Xfanout270 _07866_ vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__buf_2
Xfanout281 net283 vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__clkbuf_2
Xfanout1279 net1281 vssd1 vssd1 vccd1 vccd1 net1279 sky130_fd_sc_hd__clkbuf_4
X_16731_ clknet_leaf_69_wb_clk_i _02418_ _00714_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout292 net293 vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__clkbuf_2
X_13943_ _04218_ _04234_ vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__nor2_4
XFILLER_0_89_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16662_ clknet_leaf_12_wb_clk_i _02349_ _00645_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13874_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[8\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[9\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[10\] vssd1 vssd1 vccd1 vccd1 _04185_
+ sky130_fd_sc_hd__and3_1
X_15613_ net1240 vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__inv_2
X_12825_ net1732 net641 net609 _03646_ vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__a22o_1
X_16593_ clknet_leaf_114_wb_clk_i _02280_ _00576_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15544_ net1215 vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__inv_2
X_12756_ net363 _03597_ _03598_ net1060 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__a32o_1
XANTENNA__08607__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_7__f_wb_clk_i_X clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08834__C net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11707_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\]
+ _07800_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] vssd1 vssd1 vccd1 vccd1
+ _07903_ sky130_fd_sc_hd__a31o_1
X_15475_ net1419 vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__inv_2
XANTENNA__12129__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12687_ _07791_ _07942_ net574 vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__and3_4
XFILLER_0_25_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17214_ clknet_leaf_81_wb_clk_i _02901_ _01197_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12909__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14426_ net1308 vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__inv_2
X_11638_ net714 _07600_ vssd1 vssd1 vccd1 vccd1 _07848_ sky130_fd_sc_hd__nand2_1
XANTENNA__09235__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12924__Y _03692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10157__B _04970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11968__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08589__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17145_ clknet_leaf_102_wb_clk_i _02832_ _01128_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13582__A2 _07541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14357_ net1333 vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11569_ net3122 net153 team_01_WB.instance_to_wrap.cpu.K0.next_state vssd1 vssd1
+ vccd1 vccd1 _03272_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10396__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13319__C1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12790__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold707 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2242 sky130_fd_sc_hd__dlygate4sd3_1
X_13308_ net610 _07707_ team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1
+ vccd1 _03790_ sky130_fd_sc_hd__a21o_1
Xhold718 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2253 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_94_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold729 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2264 sky130_fd_sc_hd__dlygate4sd3_1
X_17076_ clknet_leaf_21_wb_clk_i _02763_ _01059_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14288_ net1343 vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__inv_2
XANTENNA__09665__C net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16027_ net1309 vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__inv_2
XANTENNA__12886__B1_N net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11269__A net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13239_ net2701 net354 net350 team_01_WB.instance_to_wrap.cpu.f0.i\[11\] vssd1 vssd1
+ vccd1 vccd1 _01911_ sky130_fd_sc_hd__a22o_1
X_17964__1479 vssd1 vssd1 vccd1 vccd1 _17964__1479/HI net1479 sky130_fd_sc_hd__conb_1
XANTENNA__10148__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08761__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08780_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[0\] net658 _05117_ _05118_
+ _05119_ vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__a2111o_1
Xhold1407 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2942 sky130_fd_sc_hd__dlygate4sd3_1
X_17978_ net1493 vssd1 vssd1 vccd1 vccd1 la_data_out[20] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1418 _02121_ vssd1 vssd1 vccd1 vccd1 net2953 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1429 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2964 sky130_fd_sc_hd__dlygate4sd3_1
X_16929_ clknet_leaf_54_wb_clk_i _02616_ _00912_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16568__Q team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08297__B net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10856__A0 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14047__B1 _04244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire506_X net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09401_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[27\] net699 net696 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__a22o_1
XANTENNA__10871__A3 _06065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09332_ _05665_ _05667_ _05669_ _05671_ vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__or4_1
XANTENNA__13270__A1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08744__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11281__B1 _07620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09263_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[20\] net690 net663 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_138_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout233_A net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12039__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08214_ net2418 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[59\] net1055 vssd1 vssd1
+ vccd1 vccd1 _03473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09194_ net1085 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[17\] net911
+ vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11878__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08145_ _04612_ _04613_ _04614_ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout400_A _03566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1142_A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10387__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12781__B1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08076_ _04525_ _04550_ _04551_ net569 net1564 vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_112_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15874__A net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10139__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1407_A net1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout390_X net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout488_X net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout867_A net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13394__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[6\] vssd1 vssd1 vccd1 vccd1
+ net1547 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[5\] vssd1 vssd1 vccd1 vccd1
+ net1558 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13089__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12502__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08978_ net1007 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[8\] net939 vssd1
+ vssd1 vccd1 vccd1 _05318_ sky130_fd_sc_hd__and3_1
Xhold34 team_01_WB.instance_to_wrap.a1.ADR_I\[4\] vssd1 vssd1 vccd1 vccd1 net1569
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 _01982_ vssd1 vssd1 vccd1 vccd1 net1580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 team_01_WB.instance_to_wrap.cpu.f0.write_data\[11\] vssd1 vssd1 vccd1 vccd1
+ net1591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 team_01_WB.instance_to_wrap.cpu.f0.write_data\[22\] vssd1 vssd1 vccd1 vccd1
+ net1602 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11639__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold78 net112 vssd1 vssd1 vccd1 vccd1 net1613 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[3\] vssd1 vssd1 vccd1 vccd1
+ net1624 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout655_X net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1397_X net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08504__A2 _04837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10940_ _07059_ _07061_ net517 vssd1 vssd1 vccd1 vccd1 _07280_ sky130_fd_sc_hd__mux2_1
XANTENNA__10311__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout822_X net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10871_ _05963_ _05996_ _06032_ _06065_ net548 net536 vssd1 vssd1 vccd1 vccd1 _07211_
+ sky130_fd_sc_hd__mux4_1
X_12610_ net2768 net251 net398 vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08268__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13590_ net186 _04033_ _04034_ net724 vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__a211o_1
XFILLER_0_94_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08654__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12541_ net2681 net254 net406 vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15260_ net1246 vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12472_ net2447 net261 net411 vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11788__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14211_ net2566 vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11423_ _07701_ _07702_ _07735_ net324 vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15191_ net1213 vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10378__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_9 _03654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11354_ net1070 net1071 vssd1 vssd1 vccd1 vccd1 _07683_ sky130_fd_sc_hd__nand2_1
X_14142_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[55\] _04236_ _04265_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__a22o_1
XANTENNA__10705__B net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10305_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[18\] net819 net791 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06645_ sky130_fd_sc_hd__a22o_1
XANTENNA__08991__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11285_ _07554_ _07566_ _07624_ vssd1 vssd1 vccd1 vccd1 _07625_ sky130_fd_sc_hd__or3_1
X_14073_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[68\] _04233_ _04262_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[52\]
+ vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10236_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[9\] net786 net756 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[9\]
+ _06569_ vssd1 vssd1 vccd1 vccd1 _06576_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_5_Left_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13024_ net2918 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[70\] net854 vssd1 vssd1
+ vccd1 vccd1 _02101_ sky130_fd_sc_hd__mux2_1
X_17901_ net1436 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
Xfanout1010 net1014 vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__buf_2
Xfanout1021 net1030 vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__clkbuf_2
X_17832_ clknet_leaf_120_wb_clk_i _03508_ _01772_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12412__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10167_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[10\] _04667_ net774
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[10\] vssd1 vssd1 vccd1 vccd1
+ _06507_ sky130_fd_sc_hd__a22o_1
Xfanout1032 net1033 vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__clkbuf_4
Xfanout1043 net1059 vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__buf_2
Xfanout1054 net1055 vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__clkbuf_4
Xfanout1065 team_01_WB.instance_to_wrap.cpu.RU0.state\[4\] vssd1 vssd1 vccd1 vccd1
+ net1065 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08829__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17763_ clknet_leaf_93_wb_clk_i net2322 _01703_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[33\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1076 team_01_WB.instance_to_wrap.cpu.IM0.pc_enable vssd1 vssd1 vccd1 vccd1
+ net1076 sky130_fd_sc_hd__buf_2
Xfanout1087 net1088 vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12827__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10098_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] net625 _06436_ _06437_
+ vssd1 vssd1 vccd1 vccd1 _06438_ sky130_fd_sc_hd__a22o_4
X_14975_ net1312 vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__inv_2
Xfanout1098 net1103 vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_107_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16714_ clknet_leaf_32_wb_clk_i _02401_ _00697_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13926_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__nand2b_4
XANTENNA__14029__B1 _04259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17694_ clknet_leaf_137_wb_clk_i _03378_ _01635_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_92_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10302__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16645_ clknet_leaf_52_wb_clk_i _02332_ _00628_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13857_ net1180 net1067 net2055 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[18\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_9_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12808_ net1038 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[7\] vssd1 vssd1 vccd1
+ vccd1 _03634_ sky130_fd_sc_hd__or2_2
XFILLER_0_69_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16576_ clknet_leaf_38_wb_clk_i _02263_ _00559_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09456__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13788_ _04168_ _04170_ vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__nand2_1
XANTENNA__09022__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15527_ net1391 vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_44_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12739_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] net1062 net365 _03586_
+ vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_32_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09957__A net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15458_ net1320 vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_96_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08861__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13555__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13479__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14409_ net1359 vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_133_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15389_ net1315 vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_133_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12763__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17128_ clknet_leaf_61_wb_clk_i _02815_ _01111_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold504 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2039 sky130_fd_sc_hd__dlygate4sd3_1
Xhold515 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2050 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold526 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2061 sky130_fd_sc_hd__dlygate4sd3_1
Xhold537 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2072 sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2083 sky130_fd_sc_hd__dlygate4sd3_1
Xhold559 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2094 sky130_fd_sc_hd__dlygate4sd3_1
X_09950_ net1156 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[3\] _04660_
+ vssd1 vssd1 vccd1 vccd1 _06290_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17059_ clknet_leaf_25_wb_clk_i _02746_ _01042_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_08901_ net1025 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[2\] net915 vssd1
+ vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__and3_1
X_09881_ _06165_ _06194_ _06220_ vssd1 vssd1 vccd1 vccd1 _06221_ sky130_fd_sc_hd__or3_1
XFILLER_0_148_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17682__Q team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_57_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08832_ net1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[1\] net915 vssd1
+ vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__and3_1
XANTENNA__12322__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1204 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2739 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10541__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1215 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[16\] vssd1 vssd1 vccd1 vccd1
+ net2750 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1226 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[50\] vssd1 vssd1 vccd1 vccd1
+ net2761 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08739__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1237 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[106\] vssd1 vssd1 vccd1 vccd1
+ net2772 sky130_fd_sc_hd__dlygate4sd3_1
X_08763_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[4\] net649 _05081_ _05085_
+ _05087_ vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__a2111o_1
Xhold1248 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2783 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1259 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[80\] vssd1 vssd1 vccd1 vccd1
+ net2794 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08694_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[7\] net698 _05019_ _05022_
+ _05029_ vssd1 vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_68_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1092_A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout448_A _07958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09447__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10057__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08474__C net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09315_ net1121 net711 net594 vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09998__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout615_A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout236_X net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09246_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[21\] net680 net655 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08771__A _04708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09177_ net1091 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[16\] net887
+ vssd1 vssd1 vccd1 vccd1 _05517_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout403_X net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1145_X net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08128_ _04484_ team_01_WB.instance_to_wrap.cpu.f0.num\[9\] team_01_WB.instance_to_wrap.cpu.f0.num\[12\]
+ _04482_ vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout984_A _04629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08059_ _04514_ _04528_ _04529_ _04522_ vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__o22ai_1
XANTENNA__11309__A1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11070_ _05006_ _06526_ _07374_ net340 _04969_ vssd1 vssd1 vccd1 vccd1 _07410_ sky130_fd_sc_hd__o32a_1
XANTENNA__13836__B net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout772_X net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__buf_2
XFILLER_0_101_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10021_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[1\] net798 net792 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06361_ sky130_fd_sc_hd__a22o_1
XANTENNA__08725__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12232__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10532__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08649__C net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12809__A1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12809__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14760_ net1375 vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__inv_2
XANTENNA__09686__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13482__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11972_ net1920 net238 net471 vssd1 vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__mux2_1
XANTENNA__13482__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09150__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13711_ team_01_WB.instance_to_wrap.cpu.c0.count\[15\] _04502_ _04109_ _04125_ vssd1
+ vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[16\] sky130_fd_sc_hd__a31o_1
XANTENNA__10296__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10923_ _07212_ _07256_ net525 vssd1 vssd1 vccd1 vccd1 _07263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10687__S net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14691_ net1195 vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16430_ clknet_leaf_130_wb_clk_i _02184_ _00413_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13642_ net199 net195 _07799_ _07920_ net645 vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__o2111a_1
X_10854_ net376 _06496_ vssd1 vssd1 vccd1 vccd1 _07194_ sky130_fd_sc_hd__nor2_1
XFILLER_0_156_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13234__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_39_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17963__1478 vssd1 vssd1 vccd1 vccd1 _17963__1478/HI net1478 sky130_fd_sc_hd__conb_1
XFILLER_0_27_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15779__A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16361_ clknet_leaf_99_wb_clk_i _02115_ _00344_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[84\]
+ sky130_fd_sc_hd__dfstp_1
X_13573_ _03918_ _04019_ vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__xor2_1
XFILLER_0_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10785_ net505 net333 net331 vssd1 vssd1 vccd1 vccd1 _07125_ sky130_fd_sc_hd__a21o_1
XANTENNA__11796__A1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10419__C net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15312_ net1271 vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__inv_2
X_12524_ net2289 net221 net403 vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__mux2_1
X_16292_ clknet_leaf_121_wb_clk_i _02046_ _00275_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12915__B net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15243_ net1397 vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12455_ net2364 net290 net416 vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_969 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09496__B _05835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12407__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12745__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11406_ net1069 _07694_ net323 vssd1 vssd1 vccd1 vccd1 _07726_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_62_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15174_ net1383 vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__inv_2
X_12386_ net2449 net308 net426 vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14125_ _04405_ _04406_ _04408_ _04410_ vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__or4_1
XFILLER_0_104_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11337_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[0\] team_01_WB.instance_to_wrap.cpu.f0.state\[4\]
+ _04561_ _07652_ vssd1 vssd1 vccd1 vccd1 _07667_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_150_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_150_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_123_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14056_ _04226_ _04250_ _04255_ _04264_ vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__or4_1
X_11268_ _06915_ _07365_ _07366_ net335 _07607_ vssd1 vssd1 vccd1 vccd1 _07608_ sky130_fd_sc_hd__o221a_1
XFILLER_0_120_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13007_ net2718 net2568 net856 vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__mux2_1
X_10219_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[8\] net815 net769 _06557_
+ _06558_ vssd1 vssd1 vccd1 vccd1 _06559_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12142__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11199_ net515 _07063_ _07099_ _07538_ vssd1 vssd1 vccd1 vccd1 _07539_ sky130_fd_sc_hd__a31o_1
X_17815_ clknet_leaf_100_wb_clk_i _03491_ _01755_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[85\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_89_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_89_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11981__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17746_ clknet_leaf_123_wb_clk_i net2573 _01686_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_14958_ net1298 vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09141__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13909_ _04207_ net571 _04206_ vssd1 vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_85_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17677_ clknet_leaf_157_wb_clk_i _03362_ _01618_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14889_ net1295 vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11282__A _07088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16628_ clknet_leaf_66_wb_clk_i _02315_ _00611_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09429__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13225__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16559_ clknet_leaf_0_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[25\]
+ _00542_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_135_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09100_ net1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[13\] net901
+ vssd1 vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__and3_1
XFILLER_0_128_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09031_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[9\] net700 _05348_ _05358_
+ net707 vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_26_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16581__Q team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[13\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13528__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10185__X _06525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12317__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12736__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11539__B2 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold301 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1836 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_68_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold312 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1847 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_27_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_40_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold323 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[9\] vssd1 vssd1 vccd1 vccd1
+ net1869 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08955__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold345 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1880 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 team_01_WB.instance_to_wrap.a1.ADR_I\[5\] vssd1 vssd1 vccd1 vccd1 net1891
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1902 sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1913 sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[4\] net758 net749 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06273_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold389 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[20\] vssd1 vssd1 vccd1 vccd1
+ net1924 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout803 _04643_ vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__clkbuf_4
Xfanout814 _04637_ vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__buf_4
Xfanout825 _04579_ vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__buf_2
XANTENNA_fanout398_A _03567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13161__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout836 _03737_ vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__buf_2
X_09864_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[12\] net802 net737 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06204_ sky130_fd_sc_hd__a22o_1
XANTENNA__12052__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout847 net851 vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__clkbuf_4
Xfanout858 net868 vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1105_A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout869 net873 vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11711__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10514__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1001 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2536 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1012 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2547 sky130_fd_sc_hd__dlygate4sd3_1
X_08815_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[1\] net703 vssd1 vssd1
+ vccd1 vccd1 _05155_ sky130_fd_sc_hd__or2_1
XANTENNA__09380__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08469__C net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13943__Y _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1023 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1034 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[26\] vssd1 vssd1 vccd1 vccd1
+ net2569 sky130_fd_sc_hd__dlygate4sd3_1
X_09795_ _06134_ vssd1 vssd1 vccd1 vccd1 _06135_ sky130_fd_sc_hd__inv_2
XANTENNA__11891__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1045 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2580 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout565_A net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout186_X net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1056 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[23\] vssd1 vssd1 vccd1 vccd1
+ net2591 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1067 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[39\] vssd1 vssd1 vccd1 vccd1
+ net2602 sky130_fd_sc_hd__dlygate4sd3_1
X_08746_ net1014 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[4\] net891 vssd1
+ vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_107_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1078 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2613 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_77_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1089 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2624 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13391__B _05705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08677_ net1008 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[7\] net904 vssd1
+ vssd1 vccd1 vccd1 _05017_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout732_A net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10817__A3 _06811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08485__B net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout520_X net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_66_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_9_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10570_ _04736_ _04738_ vssd1 vssd1 vccd1 vccd1 _06910_ sky130_fd_sc_hd__nand2b_2
XANTENNA__09597__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09840__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08932__C net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09229_ _04884_ _04919_ _05567_ vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__nor3_1
XANTENNA__12227__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_86_Left_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12240_ net2344 net266 net439 vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout987_X net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13858__A_N net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12171_ net2067 net234 net447 vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08800__D1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12751__A net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11122_ net370 _07386_ _07388_ net337 _07461_ vssd1 vssd1 vccd1 vccd1 _07462_ sky130_fd_sc_hd__a221o_1
Xhold890 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2425 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13152__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13058__S net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11053_ _07388_ _06340_ net518 vssd1 vssd1 vccd1 vccd1 _07393_ sky130_fd_sc_hd__and3b_1
X_15930_ net1353 vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10505__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10004_ net1156 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[1\] net953 vssd1
+ vssd1 vccd1 vccd1 _06344_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09371__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11086__B net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15861_ net1357 vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_95_Left_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17600_ clknet_leaf_86_wb_clk_i _03287_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_14812_ net1247 vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__inv_2
X_15792_ net1205 vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__inv_2
X_17531_ clknet_leaf_75_wb_clk_i _03218_ _01514_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1590 net148 vssd1 vssd1 vccd1 vccd1 net3125 sky130_fd_sc_hd__dlygate4sd3_1
X_14743_ net1197 vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__inv_2
XANTENNA__11466__B1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11955_ net2938 net318 net478 vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10906_ _04884_ _06671_ _07244_ _07245_ vssd1 vssd1 vccd1 vccd1 _07246_ sky130_fd_sc_hd__o22a_1
X_17462_ clknet_leaf_24_wb_clk_i _03149_ _01445_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14674_ net1306 vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__inv_2
XANTENNA__08882__A1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11886_ net2124 net292 net486 vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__mux2_1
X_16413_ clknet_leaf_124_wb_clk_i _02167_ _00396_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11218__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13625_ _03892_ _04063_ vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__xnor2_1
X_10837_ net334 _07176_ vssd1 vssd1 vccd1 vccd1 _07177_ sky130_fd_sc_hd__nand2_1
X_17393_ clknet_leaf_116_wb_clk_i _03080_ _01376_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09003__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09426__A3 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16344_ clknet_leaf_95_wb_clk_i _02098_ _00327_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[67\]
+ sky130_fd_sc_hd__dfrtp_1
X_13556_ _03923_ _03924_ vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__nor2_1
XANTENNA__09831__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10768_ _06314_ _07055_ vssd1 vssd1 vccd1 vccd1 _07108_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12507_ net2137 net257 net409 vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__mux2_1
X_16275_ clknet_leaf_88_wb_clk_i _00003_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[4\]
+ sky130_fd_sc_hd__dfxtp_4
XANTENNA__12137__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13487_ _03845_ _03946_ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10699_ _06948_ _06953_ net535 vssd1 vssd1 vccd1 vccd1 _07039_ sky130_fd_sc_hd__mux2_1
X_18014_ net636 vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_130_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15226_ net1371 vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12438_ net2506 net267 net415 vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11976__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15157_ net1282 vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12369_ net2312 net269 net423 vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__mux2_1
X_14108_ _04385_ _04394_ vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09673__C net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15088_ net1273 vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14039_ net1568 net605 _04328_ net1183 vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_56_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09362__A2 _04766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13763__Y _04152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14588__A net1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08600_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[15\] net689 _04923_
+ _04925_ _04926_ vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__a2111o_1
X_09580_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[25\] net788 net757 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[25\]
+ _05919_ vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__a221o_1
XANTENNA__12600__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08586__A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16576__Q team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08531_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[18\] net654 _04850_
+ _04855_ _04868_ vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__a2111o_1
X_17729_ clknet_leaf_136_wb_clk_i team_01_WB.instance_to_wrap.cpu.f0.next_write_i
+ _01669_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_i sky130_fd_sc_hd__dfrtp_4
XANTENNA__13997__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_100_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_77_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08462_ net1001 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[23\] net925 vssd1
+ vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_102_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08393_ _04709_ _04732_ vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_154_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10125__A1_N net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08752__C net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_150_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12047__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1055_A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09014_ net1021 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[9\] net927 vssd1
+ vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__and3_1
XANTENNA__13938__Y _04230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11886__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold120 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 net1655
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold131 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[12\] vssd1 vssd1 vccd1 vccd1
+ net1666 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[10\] vssd1 vssd1 vccd1 vccd1
+ net1677 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1222_A net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10735__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold153 team_01_WB.instance_to_wrap.cpu.f0.write_data\[25\] vssd1 vssd1 vccd1 vccd1
+ net1688 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold164 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[7\] vssd1 vssd1 vccd1 vccd1
+ net1699 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[23\] vssd1 vssd1 vccd1 vccd1
+ net1710 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout682_A net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold186 _03340_ vssd1 vssd1 vccd1 vccd1 net1721 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout600 _04754_ vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10803__B net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold197 team_01_WB.instance_to_wrap.a1.ADR_I\[3\] vssd1 vssd1 vccd1 vccd1 net1732
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout611 net614 vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11187__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13134__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13954__X _04246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17962__1477 vssd1 vssd1 vccd1 vccd1 _17962__1477/HI net1477 sky130_fd_sc_hd__conb_1
X_09916_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[4\] net752 net742 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06256_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout622 net623 vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1010_X net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout633 _03733_ vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__clkbuf_4
Xfanout644 _04839_ vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10522__C net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout655 _04817_ vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__buf_4
Xfanout666 _04804_ vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__buf_4
XANTENNA__09353__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11696__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09847_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[13\] net763 net622 vssd1
+ vssd1 vccd1 vccd1 _06187_ sky130_fd_sc_hd__o21a_1
Xfanout677 _04790_ vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__buf_2
Xfanout688 _04773_ vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_126_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout470_X net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout699 _04760_ vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_126_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout568_X net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12510__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13437__A1 team_01_WB.instance_to_wrap.cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09778_ _06113_ _06114_ _06115_ _06117_ vssd1 vssd1 vccd1 vccd1 _06118_ sky130_fd_sc_hd__or4_1
XANTENNA__08927__C net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09105__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08729_ _05065_ _05066_ _05067_ _05068_ vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__or4_1
XANTENNA__13988__A2 _04241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_723 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout735_X net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11740_ _07797_ _07929_ vssd1 vssd1 vccd1 vccd1 _07930_ sky130_fd_sc_hd__nor2_1
XANTENNA__10120__B1 _04667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout902_X net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11671_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[17\] _07232_ net713 vssd1 vssd1
+ vccd1 vccd1 _07874_ sky130_fd_sc_hd__mux2_1
X_13410_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] _05220_ vssd1 vssd1 vccd1
+ vccd1 _03871_ sky130_fd_sc_hd__or2_1
X_10622_ _05839_ _06826_ _06828_ vssd1 vssd1 vccd1 vccd1 _06962_ sky130_fd_sc_hd__nand3_1
XFILLER_0_10_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14390_ net1193 vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__inv_2
X_13341_ _07681_ _03815_ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10553_ _06891_ _06892_ net538 vssd1 vssd1 vccd1 vccd1 _06893_ sky130_fd_sc_hd__mux2_1
XANTENNA__08007__Y _04504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10974__A2 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16060_ clknet_leaf_154_wb_clk_i _01853_ _00048_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\]
+ sky130_fd_sc_hd__dfrtp_4
X_13272_ net1068 _03748_ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10484_ _06750_ _06819_ _06823_ vssd1 vssd1 vccd1 vccd1 _06824_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11796__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15011_ net1250 vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__inv_2
X_12223_ _07790_ _07791_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[11\] vssd1 vssd1
+ vccd1 vccd1 _07960_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09041__A1 net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12154_ net2295 net317 net454 vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13125__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15792__A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11105_ _07282_ _07285_ net516 vssd1 vssd1 vccd1 vccd1 _07445_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16962_ clknet_leaf_55_wb_clk_i _02649_ _00945_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12085_ net2534 net293 net462 vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__mux2_1
XANTENNA__13676__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11036_ _05006_ _06527_ vssd1 vssd1 vccd1 vccd1 _07376_ sky130_fd_sc_hd__or2_1
X_15913_ net1402 vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__inv_2
X_16893_ clknet_leaf_66_wb_clk_i _02580_ _00876_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15844_ net1325 vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__inv_2
XANTENNA__12420__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15775_ net1199 vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__inv_2
XANTENNA__13979__A2 _04221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12987_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[99\] net2532 net862 vssd1 vssd1
+ vccd1 vccd1 _02138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09789__X _06129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14726_ net1209 vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__inv_2
X_17514_ clknet_leaf_10_wb_clk_i _03201_ _01497_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10111__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11938_ net2278 net239 net475 vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17445_ clknet_leaf_51_wb_clk_i _03132_ _01428_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10662__A1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14657_ net1218 vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11869_ net2995 net200 net484 vssd1 vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__mux2_1
XANTENNA__13104__X _03728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13608_ net720 _07520_ net1073 vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__o21a_1
XANTENNA__15032__A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17376_ clknet_leaf_47_wb_clk_i _03063_ _01359_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09804__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14588_ net1408 vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__inv_2
XANTENNA__09668__C net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16327_ clknet_leaf_91_wb_clk_i _02081_ _00310_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[50\]
+ sky130_fd_sc_hd__dfrtp_1
X_13539_ _03928_ _03931_ _03990_ _03927_ vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_31_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08083__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_859 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16258_ clknet_leaf_156_wb_clk_i net1736 _00246_ vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15209_ net1288 vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10178__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16189_ clknet_leaf_1_wb_clk_i _01949_ _00177_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10904__A net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09583__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13116__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10342__C net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09701_ net1154 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[21\] net985
+ vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__and3_1
XANTENNA__09335__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17690__Q team_01_WB.instance_to_wrap.cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11142__A2 _06903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11294__X _07634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09632_ net1135 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[23\] net970
+ vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_143_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12330__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08747__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09563_ net997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[25\] net952 vssd1
+ vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout263_A _07880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08514_ net1001 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[18\] net918 vssd1
+ vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__and3_1
X_09494_ team_01_WB.instance_to_wrap.cpu.CU0.bit30 net710 net594 vssd1 vssd1 vccd1
+ vccd1 _05834_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10653__A1 _04706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08445_ net1122 net1125 net1117 net1120 vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__and4bb_4
XANTENNA_fanout430_A _07965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1172_A team_01_WB.instance_to_wrap.cpu.DM0.ihit vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_18_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout528_A net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08376_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] _04715_ _04710_ vssd1 vssd1
+ vccd1 vccd1 _04716_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08482__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1058_X net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14147__A2 _04221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout897_A _04793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12505__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10169__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11188__Y _07528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout685_X net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1406 net1408 vssd1 vssd1 vccd1 vccd1 net1406 sky130_fd_sc_hd__buf_4
Xfanout1417 net1418 vssd1 vssd1 vccd1 vccd1 net1417 sky130_fd_sc_hd__buf_4
XANTENNA__11118__C1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11348__C net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13658__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1428 net1429 vssd1 vssd1 vccd1 vccd1 net1428 sky130_fd_sc_hd__clkbuf_4
Xfanout430 _07965_ vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__clkbuf_4
Xfanout441 _07962_ vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__buf_6
Xfanout452 _07957_ vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__buf_4
XANTENNA__09326__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout463 _07954_ vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_6_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout474 _07952_ vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11133__A2 _06924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout485 _07948_ vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__buf_6
X_12910_ _04918_ net577 net360 vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__o21ba_1
Xfanout496 net498 vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__buf_6
XANTENNA__12240__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13890_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[0\] net572 vssd1 vssd1 vccd1
+ vccd1 _03247_ sky130_fd_sc_hd__and2b_1
XANTENNA__10892__A1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12841_ net2027 net273 net380 vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15560_ net1398 vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__inv_2
X_12772_ net1895 net639 net607 _03609_ vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14511_ net1400 vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__inv_2
X_11723_ _07800_ _07915_ vssd1 vssd1 vccd1 vccd1 _07916_ sky130_fd_sc_hd__nor2_1
X_15491_ net1270 vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11380__A team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_7_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17230_ clknet_leaf_28_wb_clk_i _02917_ _01213_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_14442_ net1227 vssd1 vssd1 vccd1 vccd1 _00236_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11654_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] _07814_ vssd1 vssd1
+ vccd1 vccd1 _07861_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17161_ clknet_leaf_40_wb_clk_i _02848_ _01144_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10605_ _06938_ _06944_ net519 vssd1 vssd1 vccd1 vccd1 _06945_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14373_ net1208 vssd1 vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11585_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] _07801_ vssd1 vssd1 vccd1
+ vccd1 _07802_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16112_ clknet_leaf_138_wb_clk_i _01887_ _00100_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13324_ team_01_WB.instance_to_wrap.cpu.f0.i\[17\] _07703_ vssd1 vssd1 vccd1 vccd1
+ _03803_ sky130_fd_sc_hd__nor2_1
XANTENNA__14138__A2 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17092_ clknet_leaf_82_wb_clk_i _02779_ _01075_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10536_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[31\] net664 net650 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06876_ sky130_fd_sc_hd__a22o_1
Xwire886 _04803_ vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__clkbuf_2
X_16043_ clknet_leaf_88_wb_clk_i _01837_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13255_ team_01_WB.instance_to_wrap.cpu.f0.i\[25\] team_01_WB.instance_to_wrap.cpu.f0.i\[24\]
+ _03746_ vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__and3_1
XANTENNA__12415__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10467_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[26\] net783 _06786_ _06788_
+ _06793_ vssd1 vssd1 vccd1 vccd1 _06807_ sky130_fd_sc_hd__a2111o_1
X_12206_ net2626 net262 net444 vssd1 vssd1 vccd1 vccd1 _02783_ sky130_fd_sc_hd__mux2_1
XANTENNA__11098__Y _07438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_57_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13186_ net23 net835 net628 net1724 vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__o22a_1
X_10398_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] _06737_ net623 vssd1
+ vssd1 vccd1 vccd1 _06738_ sky130_fd_sc_hd__mux2_2
X_12137_ net1809 net237 net451 vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__mux2_1
XANTENNA__13649__A1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17994_ net635 vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09317__A2 _05654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16945_ clknet_leaf_113_wb_clk_i _02632_ _00928_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_12068_ net1827 net200 net459 vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__mux2_1
XANTENNA__09951__C net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08848__B _05153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12150__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11019_ _07127_ _07358_ vssd1 vssd1 vccd1 vccd1 _07359_ sky130_fd_sc_hd__nand2_1
X_16876_ clknet_leaf_20_wb_clk_i _02563_ _00859_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08567__C net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15827_ net1338 vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__inv_2
XANTENNA__12938__X _03702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15758_ net1341 vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_32_Left_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14709_ net1193 vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__inv_2
X_15689_ net1295 vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11290__A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08230_ net2694 net2482 net1054 vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__mux2_1
X_17428_ clknet_leaf_66_wb_clk_i _03115_ _01411_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_17961__1476 vssd1 vssd1 vccd1 vccd1 _17961__1476/HI net1476 sky130_fd_sc_hd__conb_1
XFILLER_0_28_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08161_ net1757 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[112\] net1047 vssd1 vssd1
+ vccd1 vccd1 _03526_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17359_ clknet_leaf_31_wb_clk_i _03046_ _01342_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09695__A net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08092_ team_01_WB.instance_to_wrap.cpu.K0.keyvalid _04531_ vssd1 vssd1 vccd1 vccd1
+ _04563_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17685__Q team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_42_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload40 clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload40/Y sky130_fd_sc_hd__inv_6
Xclkload51 clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload51/Y sky130_fd_sc_hd__inv_8
XPHY_EDGE_ROW_41_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12325__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload62 clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload62/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload73 clknet_leaf_56_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload73/Y sky130_fd_sc_hd__inv_6
XFILLER_0_141_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload84 clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload84/X sky130_fd_sc_hd__clkbuf_8
Xclkload95 clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload95/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_114_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08994_ net1087 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[8\] net900 vssd1
+ vssd1 vccd1 vccd1 _05334_ sky130_fd_sc_hd__and3_1
XANTENNA__10072__C net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1018_A net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout380_A net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12312__A1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout478_A _07950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12060__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09615_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[24\] net746 _05938_ _05941_
+ _05944_ vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13951__Y _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10874__A1 _06779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11752__X _07939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1387_A net1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09546_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[28\] net805 net731 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout812_A net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09477_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[30\] net672 net658 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout433_X net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1175_X net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08428_ net1108 net927 vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__and2_1
XFILLER_0_109_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13576__B1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload1 clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload1/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__09101__C net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout600_X net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08047__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08359_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[30\] net739 _04668_ _04664_
+ _04655_ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_46_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11370_ net324 vssd1 vssd1 vccd1 vccd1 _07699_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08940__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10321_ net990 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[18\] net984 vssd1
+ vssd1 vccd1 vccd1 _06661_ sky130_fd_sc_hd__and3_1
XANTENNA__12235__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13040_ net2687 net2629 net854 vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__mux2_1
XANTENNA__09547__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10252_ net560 _05338_ _06564_ vssd1 vssd1 vccd1 vccd1 _06592_ sky130_fd_sc_hd__o21ba_1
X_10183_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[10\] _04678_ _06522_
+ vssd1 vssd1 vccd1 vccd1 _06523_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10831__X _07171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1203 net1205 vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__buf_4
Xfanout1214 net1216 vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1225 net1226 vssd1 vssd1 vccd1 vccd1 net1225 sky130_fd_sc_hd__buf_4
Xfanout1236 net1237 vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__buf_4
X_14991_ net1295 vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__inv_2
Xfanout1247 net1248 vssd1 vssd1 vccd1 vccd1 net1247 sky130_fd_sc_hd__buf_4
XANTENNA_input39_A wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1258 net1269 vssd1 vssd1 vccd1 vccd1 net1258 sky130_fd_sc_hd__buf_4
Xfanout260 _07888_ vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__buf_1
Xfanout1269 net1303 vssd1 vssd1 vccd1 vccd1 net1269 sky130_fd_sc_hd__clkbuf_4
Xfanout271 _07866_ vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__buf_2
Xfanout282 net283 vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__buf_2
X_16730_ clknet_leaf_78_wb_clk_i _02417_ _00713_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09116__Y _05456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13942_ _04222_ _04228_ vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__nand2_2
Xfanout293 net295 vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08020__Y _04516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10865__A1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16661_ clknet_leaf_115_wb_clk_i _02348_ _00644_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13873_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[4\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[7\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__or4_1
XANTENNA__10865__B2 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15612_ net1245 vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__inv_2
X_12824_ net364 _03644_ _03645_ net1063 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__a32o_1
X_16592_ clknet_leaf_148_wb_clk_i _02279_ _00575_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_104_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_104_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15543_ net1215 vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__inv_2
X_12755_ net1034 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[24\] vssd1 vssd1 vccd1
+ vccd1 _03598_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10093__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11706_ net718 _07531_ net616 _07901_ vssd1 vssd1 vccd1 vccd1 _07902_ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15474_ net1286 vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__inv_2
X_12686_ net1777 net289 net388 vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17213_ clknet_leaf_65_wb_clk_i _02900_ _01196_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_14425_ net1342 vssd1 vssd1 vccd1 vccd1 _00219_ sky130_fd_sc_hd__inv_2
X_11637_ net1957 net206 net501 vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09011__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17144_ clknet_leaf_49_wb_clk_i _02831_ _01127_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14356_ net1333 vssd1 vssd1 vccd1 vccd1 _00150_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_42_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11568_ team_01_WB.instance_to_wrap.cpu.K0.count\[1\] team_01_WB.instance_to_wrap.cpu.K0.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__nand2b_1
XANTENNA__09946__C net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13307_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[23\] net826 _03787_ _03789_
+ vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__o22a_1
XANTENNA__12790__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold708 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2243 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold719 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2254 sky130_fd_sc_hd__dlygate4sd3_1
X_10519_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[31\] net695 net661 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06859_ sky130_fd_sc_hd__a22o_1
X_17075_ clknet_leaf_22_wb_clk_i _02762_ _01058_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14287_ net1337 vssd1 vssd1 vccd1 vccd1 _00081_ sky130_fd_sc_hd__inv_2
XANTENNA__10454__A net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12145__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11499_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[13\] _07756_ vssd1 vssd1 vccd1
+ vccd1 _07777_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_94_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16026_ net1309 vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__inv_2
X_13238_ net2582 net354 net350 team_01_WB.instance_to_wrap.cpu.f0.i\[12\] vssd1 vssd1
+ vccd1 vccd1 _01912_ sky130_fd_sc_hd__a22o_1
XANTENNA__11984__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13169_ net137 net848 net840 net1689 vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__a22o_1
XANTENNA__08859__A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17977_ net1492 vssd1 vssd1 vccd1 vccd1 la_data_out[19] sky130_fd_sc_hd__buf_2
Xhold1408 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[106\] vssd1 vssd1 vccd1 vccd1
+ net2943 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1419 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2954 sky130_fd_sc_hd__dlygate4sd3_1
X_16928_ clknet_leaf_46_wb_clk_i _02615_ _00911_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_140_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10305__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09710__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16859_ clknet_leaf_71_wb_clk_i _02546_ _00842_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09400_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[27\] net680 net658 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_49_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09331_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[24\] net692 net648 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[24\]
+ _05670_ vssd1 vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10084__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11281__A1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09262_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[20\] net695 _05600_
+ _05601_ vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_138_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08213_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[68\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[60\]
+ net1045 vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09193_ net1005 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[17\] net925 vssd1
+ vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__and3_1
XANTENNA__09226__A1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout226_A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08144_ team_01_WB.instance_to_wrap.cpu.f0.i\[30\] _04493_ _04496_ team_01_WB.instance_to_wrap.cpu.f0.i\[6\]
+ _04590_ vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__o221a_1
XFILLER_0_16_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09777__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12781__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload140 clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload140/Y sky130_fd_sc_hd__inv_8
XFILLER_0_70_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12055__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08075_ team_01_WB.instance_to_wrap.cpu.f0.i\[4\] _04524_ vssd1 vssd1 vccd1 vccd1
+ _04551_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1135_A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout595_A net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11894__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1302_A net1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10544__B1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold13 team_01_WB.instance_to_wrap.cpu.DM0.state\[1\] vssd1 vssd1 vccd1 vccd1 net1548
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ net1008 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[8\] net904 vssd1
+ vssd1 vccd1 vccd1 _05317_ sky130_fd_sc_hd__and3_1
Xhold24 team_01_WB.instance_to_wrap.a1.ADR_I\[25\] vssd1 vssd1 vccd1 vccd1 net1559
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 _02002_ vssd1 vssd1 vccd1 vccd1 net1570 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout383_X net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold46 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[3\] vssd1 vssd1 vccd1 vccd1 net1581
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11195__A net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_2_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold57 team_01_WB.instance_to_wrap.cpu.f0.write_data\[24\] vssd1 vssd1 vccd1 vccd1
+ net1592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 net123 vssd1 vssd1 vccd1 vccd1 net1603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 _01979_ vssd1 vssd1 vccd1 vccd1 net1614 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10847__A1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout648_X net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10870_ _06098_ _06636_ _06671_ _06707_ net549 net538 vssd1 vssd1 vccd1 vccd1 _07210_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_39_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08935__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09529_ net513 _05868_ vssd1 vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__and2_1
XANTENNA__09465__A1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10098__X _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout815_X net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12540_ net2633 net257 net405 vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1062 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12471_ net3171 net266 net411 vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__mux2_1
XANTENNA__12754__A net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14210_ net3066 vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11422_ team_01_WB.instance_to_wrap.cpu.f0.i\[15\] _07689_ vssd1 vssd1 vccd1 vccd1
+ _07735_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15190_ net1253 vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09768__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08670__C net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14141_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[39\] _04230_ _04259_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[23\]
+ _04425_ vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__a221o_1
X_11353_ team_01_WB.instance_to_wrap.cpu.f0.i\[14\] team_01_WB.instance_to_wrap.cpu.f0.i\[13\]
+ _07679_ vssd1 vssd1 vccd1 vccd1 _07682_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10304_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[18\] net755 net734 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06644_ sky130_fd_sc_hd__a22o_1
X_14072_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[60\] _04258_ _04266_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[20\]
+ _04359_ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__a221o_1
X_11284_ _07135_ _07611_ _07621_ _07623_ vssd1 vssd1 vccd1 vccd1 _07624_ sky130_fd_sc_hd__or4_1
XFILLER_0_120_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17900_ net1435 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
XFILLER_0_30_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13023_ net2790 net2678 net856 vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__mux2_1
X_10235_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[9\] net817 _06573_ _06574_
+ vssd1 vssd1 vccd1 vccd1 _06575_ sky130_fd_sc_hd__a211o_1
Xfanout1000 net1003 vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__buf_1
Xfanout1011 net1013 vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__clkbuf_2
Xfanout1022 net1024 vssd1 vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__clkbuf_2
X_17831_ clknet_leaf_98_wb_clk_i _03507_ _01771_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[101\]
+ sky130_fd_sc_hd__dfstp_1
X_10166_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[10\] net747 net744 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06506_ sky130_fd_sc_hd__a22o_1
Xfanout1033 team_01_WB.instance_to_wrap.cpu.RU0.InstrRead vssd1 vssd1 vccd1 vccd1
+ net1033 sky130_fd_sc_hd__buf_2
XANTENNA__09940__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17960__1475 vssd1 vssd1 vccd1 vccd1 _17960__1475/HI net1475 sky130_fd_sc_hd__conb_1
Xfanout1044 net1045 vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__clkbuf_4
Xfanout1055 net1058 vssd1 vssd1 vccd1 vccd1 net1055 sky130_fd_sc_hd__clkbuf_2
Xfanout1066 net1067 vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__clkbuf_2
X_17762_ clknet_leaf_123_wb_clk_i _03438_ _01702_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[32\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1077 net1079 vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__buf_2
Xfanout1088 net1089 vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__clkbuf_2
X_14974_ net1316 vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__inv_2
X_10097_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[7\] net763 net622 vssd1
+ vssd1 vccd1 vccd1 _06437_ sky130_fd_sc_hd__o21a_1
Xfanout1099 net1103 vssd1 vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__buf_2
X_16713_ clknet_leaf_36_wb_clk_i _02400_ _00696_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14029__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13925_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__and2b_2
XANTENNA__10838__B2 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09006__C net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17693_ clknet_leaf_137_wb_clk_i _03377_ _01634_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[14\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_clkload4_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16644_ clknet_leaf_84_wb_clk_i _02331_ _00627_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13856_ net1180 net1067 net3183 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[17\]
+ sky130_fd_sc_hd__and3b_1
XANTENNA__09303__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12807_ net1035 _07308_ vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__nand2_1
X_16575_ clknet_leaf_39_wb_clk_i _02262_ _00558_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_13787_ _04168_ _04170_ vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__or2_1
X_10999_ _07062_ _07338_ _07337_ _07333_ vssd1 vssd1 vccd1 vccd1 _07339_ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15526_ net1382 vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_106_Left_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12738_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[29\] _07056_ net1036 vssd1 vssd1
+ vccd1 vccd1 _03586_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11979__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15457_ net1239 vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12669_ net2963 net266 net387 vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14408_ net1358 vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_72_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15388_ net1245 vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14339_ net1341 vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__inv_2
X_17127_ clknet_leaf_104_wb_clk_i _02814_ _01110_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold505 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2040 sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2051 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold527 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2073 sky130_fd_sc_hd__dlygate4sd3_1
X_17058_ clknet_leaf_76_wb_clk_i _02745_ _01041_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold549 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2084 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08900_ net1107 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[2\] net942 vssd1
+ vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__and3_1
X_16009_ net1357 vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_115_Left_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12603__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10471__X _06811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09880_ _06218_ _06219_ vssd1 vssd1 vccd1 vccd1 _06220_ sky130_fd_sc_hd__nand2_1
XANTENNA__10526__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09392__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08831_ net1022 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[1\] net899 vssd1
+ vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__and3_1
XANTENNA__09931__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10631__B _06857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1205 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1216 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2751 sky130_fd_sc_hd__dlygate4sd3_1
X_08762_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[4\] net674 _05086_ _05093_
+ _05099_ vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__a2111o_1
Xhold1227 _03464_ vssd1 vssd1 vccd1 vccd1 net2762 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1055 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1238 _02137_ vssd1 vssd1 vccd1 vccd1 net2773 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1249 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2784 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10350__C net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08693_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[7\] net679 _05010_ _05017_
+ _05028_ vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_68_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08755__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_124_Left_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout343_A _04748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1085_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09314_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[22\] net701 _05648_ _05653_
+ vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__o22a_4
XANTENNA_clkbuf_leaf_56_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11254__A1 _06906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11254__B2 _05263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09998__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11889__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09245_ _05578_ _05580_ _05584_ vssd1 vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout510_A _05996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout608_A _03583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08771__B net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1252_A net1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09176_ net1010 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[16\] net917 vssd1
+ vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10365__Y _06705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08127_ _04468_ team_01_WB.instance_to_wrap.cpu.f0.num\[27\] team_01_WB.instance_to_wrap.cpu.f0.num\[24\]
+ _04471_ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__o22a_1
XFILLER_0_32_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10765__A0 _04706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1040_X net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09883__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_133_Left_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08058_ net1763 net569 _04525_ _04535_ vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout598_X net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11309__A2 _07438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout977_A _04635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12513__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10517__B1 _06855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10020_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[1\] net753 net746 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06360_ sky130_fd_sc_hd__a22o_1
XANTENNA__09383__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout765_X net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout932_X net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11971_ net2882 net271 net471 vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_95_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08489__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13710_ team_01_WB.instance_to_wrap.cpu.c0.count\[16\] _04111_ _04119_ vssd1 vssd1
+ vccd1 vccd1 _04125_ sky130_fd_sc_hd__and3_1
XANTENNA__10296__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10922_ _06904_ _07261_ vssd1 vssd1 vccd1 vccd1 _07262_ sky130_fd_sc_hd__nor2_1
X_14690_ net1202 vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13641_ _03865_ _03881_ vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__xnor2_1
X_10853_ _06530_ _07191_ _06501_ vssd1 vssd1 vccd1 vccd1 _07193_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_13_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10048__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16360_ clknet_leaf_98_wb_clk_i _02114_ _00343_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[83\]
+ sky130_fd_sc_hd__dfrtp_1
X_13572_ _03857_ _03858_ vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__and2b_1
X_10784_ _06893_ _06938_ net519 vssd1 vssd1 vccd1 vccd1 _07124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15311_ net1386 vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__inv_2
XANTENNA__11799__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12523_ net2008 net190 net403 vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16291_ clknet_leaf_116_wb_clk_i _02045_ _00274_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15242_ net1374 vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12454_ net2578 net313 net417 vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11405_ team_01_WB.instance_to_wrap.cpu.f0.i\[23\] _07712_ _07713_ net326 vssd1 vssd1
+ vccd1 vccd1 _03386_ sky130_fd_sc_hd__o211a_1
X_15173_ net1286 vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_970 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12385_ net2288 net309 net424 vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input61_X net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09793__A net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14124_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[38\] _04221_ _04261_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[118\]
+ _04409_ vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__a221o_1
X_11336_ _07666_ net1872 _07655_ vssd1 vssd1 vccd1 vccd1 _03396_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14055_ _04230_ _04243_ _04249_ _04256_ vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__or4_1
X_11267_ _04948_ _07606_ vssd1 vssd1 vccd1 vccd1 _07607_ sky130_fd_sc_hd__nand2_1
XANTENNA__10508__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13006_ net2794 net2668 net868 vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__mux2_1
XANTENNA__09374__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10218_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[8\] net756 _06539_ _06540_
+ _06546_ vssd1 vssd1 vccd1 vccd1 _06558_ sky130_fd_sc_hd__a2111o_1
X_11198_ _07100_ _07280_ _07361_ _07537_ _07535_ vssd1 vssd1 vccd1 vccd1 _07538_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_37_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11181__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17814_ clknet_leaf_99_wb_clk_i _03490_ _01754_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[84\]
+ sky130_fd_sc_hd__dfstp_1
X_10149_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[11\] net754 net730 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06489_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_89_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17745_ clknet_leaf_120_wb_clk_i _03421_ _01685_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_14957_ net1265 vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__inv_2
XANTENNA__10878__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15035__A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13908_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[7\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[8\]
+ _04204_ vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__and3_1
XANTENNA__10287__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11484__B2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17676_ clknet_leaf_158_wb_clk_i _03361_ _01617_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14888_ net1387 vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__inv_2
XANTENNA__11282__B _07154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08575__C net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10692__C1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16627_ clknet_leaf_16_wb_clk_i _02314_ _00610_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13839_ net1179 net1066 net3177 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[0\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_147_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11236__A1 _06906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11236__B2 _05263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16558_ clknet_leaf_0_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[24\]
+ _00541_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15509_ net1285 vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16489_ clknet_leaf_156_wb_clk_i _02243_ _00472_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09030_ _05366_ _05367_ _05368_ _05369_ vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__or4_2
XFILLER_0_116_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold302 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[13\] vssd1 vssd1 vccd1 vccd1
+ net1837 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10345__C net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold313 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1848 sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1859 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10211__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold335 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1881 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1892 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold368 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1903 sky130_fd_sc_hd__dlygate4sd3_1
X_09932_ _06268_ _06269_ _06270_ _06271_ vssd1 vssd1 vccd1 vccd1 _06272_ sky130_fd_sc_hd__or4_1
Xhold379 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1914 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12333__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout804 _04643_ vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__buf_6
Xfanout815 net816 vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09365__B1 _04841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09208__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout826 _04579_ vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__clkbuf_2
X_09863_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[12\] net822 net762 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06203_ sky130_fd_sc_hd__a22o_1
XANTENNA__09904__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout837 _03736_ vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__buf_2
Xfanout848 net849 vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__buf_2
XANTENNA_fanout293_A net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11172__B1 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout859 net860 vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16102__Q team_01_WB.instance_to_wrap.cpu.f0.data_adr\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08814_ _04708_ net725 net718 _04838_ net1124 vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__o41a_1
XANTENNA__11711__A2 _07269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1002 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1013 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1024 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2559 sky130_fd_sc_hd__dlygate4sd3_1
X_09794_ net374 _06131_ vssd1 vssd1 vccd1 vccd1 _06134_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout1000_A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1035 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2570 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10080__C net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1046 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2581 sky130_fd_sc_hd__dlygate4sd3_1
X_08745_ net1099 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[4\] net932 vssd1
+ vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_107_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1057 _03429_ vssd1 vssd1 vccd1 vccd1 net2592 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout460_A _07955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1068 _02078_ vssd1 vssd1 vccd1 vccd1 net2603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1079 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2614 sky130_fd_sc_hd__dlygate4sd3_1
X_08676_ net1086 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[7\] net923 vssd1
+ vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_124_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_124_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout725_A net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1088_X net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12508__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout513_X net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09228_ _04970_ _05379_ _05494_ _05567_ vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__nor4_1
XFILLER_0_1_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12727__A1 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09159_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[16\] net646 _05496_
+ _05497_ _05498_ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_32_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12170_ net1741 net239 net447 vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__mux2_1
XANTENNA__13847__B team_01_WB.instance_to_wrap.cpu.RU0.state\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout882_X net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11121_ net527 _07460_ vssd1 vssd1 vccd1 vccd1 _07461_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12243__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold880 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2415 sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2426 sky130_fd_sc_hd__dlygate4sd3_1
X_11052_ net527 _06313_ vssd1 vssd1 vccd1 vccd1 _07392_ sky130_fd_sc_hd__nor2_1
X_10003_ _06340_ _06342_ vssd1 vssd1 vccd1 vccd1 _06343_ sky130_fd_sc_hd__nor2_1
X_15860_ net1349 vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__inv_2
XANTENNA_input21_A DAT_I[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14101__B1 _04258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14811_ net1254 vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__inv_2
XANTENNA__10698__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15791_ net1191 vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__inv_2
X_17904__1439 vssd1 vssd1 vccd1 vccd1 _17904__1439/HI net1439 sky130_fd_sc_hd__conb_1
Xhold1580 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net3115 sky130_fd_sc_hd__dlygate4sd3_1
X_17530_ clknet_leaf_76_wb_clk_i _03217_ _01513_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1591 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net3126 sky130_fd_sc_hd__dlygate4sd3_1
X_11954_ net2282 net306 net478 vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__mux2_1
X_14742_ net1194 vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10905_ _04884_ net331 _07243_ net333 net369 vssd1 vssd1 vccd1 vccd1 _07245_ sky130_fd_sc_hd__a221o_1
X_14673_ net1225 vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__inv_2
X_17461_ clknet_leaf_111_wb_clk_i _03148_ _01444_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11885_ net2715 net296 net486 vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08882__A2 _05219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11218__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13624_ _03893_ _04051_ vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__nand2b_1
X_16412_ clknet_leaf_124_wb_clk_i _02166_ _00395_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10836_ _05491_ _06159_ vssd1 vssd1 vccd1 vccd1 _07176_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_15_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17392_ clknet_leaf_148_wb_clk_i _03079_ _01375_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16343_ clknet_leaf_90_wb_clk_i net2595 _00326_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[66\]
+ sky130_fd_sc_hd__dfrtp_1
X_13555_ net986 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] _04004_ _04005_
+ vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12418__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10767_ net522 _07106_ _06965_ vssd1 vssd1 vccd1 vccd1 _07107_ sky130_fd_sc_hd__a21bo_1
XANTENNA__10977__A0 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12506_ net2844 net229 net409 vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__mux2_1
X_16274_ clknet_leaf_88_wb_clk_i _00002_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13486_ _03846_ _03847_ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10698_ _07036_ _07037_ net520 vssd1 vssd1 vccd1 vccd1 _07038_ sky130_fd_sc_hd__mux2_1
X_18013_ net1511 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_130_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15225_ net1237 vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_130_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12437_ net2129 net234 net415 vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09595__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15156_ net1400 vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12368_ net2191 net243 net425 vssd1 vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__mux2_1
XANTENNA__09954__C net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14107_ _04387_ _04389_ _04391_ _04393_ vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__or4_1
X_11319_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[7\] net1176 vssd1 vssd1 vccd1
+ vccd1 _07656_ sky130_fd_sc_hd__and2_1
X_15087_ net1299 vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__inv_2
XANTENNA__12153__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12299_ net2301 net274 net433 vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__mux2_1
XANTENNA__13143__A1 net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09347__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14038_ _04319_ _04325_ _04326_ _04327_ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_56_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08867__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15989_ net1416 vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08530_ net1078 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[18\] net891
+ vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__and3_1
X_17728_ clknet_leaf_93_wb_clk_i _03405_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_08461_ net1028 net927 vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__and2_2
X_17659_ clknet_leaf_4_wb_clk_i _03344_ _01600_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_102_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08873__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09698__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08392_ net1169 _04713_ net709 vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_154_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12328__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08625__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10432__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09013_ net1094 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[9\] net939 vssd1
+ vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__and3_1
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout306_A _07935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10075__C net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold110 _02000_ vssd1 vssd1 vccd1 vccd1 net1645 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09586__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold121 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[4\] vssd1 vssd1 vccd1 vccd1 net1656
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold132 _03343_ vssd1 vssd1 vccd1 vccd1 net1667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 net127 vssd1 vssd1 vccd1 vccd1 net1678 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold154 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[7\] vssd1 vssd1 vccd1 vccd1 net1689
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 team_01_WB.instance_to_wrap.cpu.f0.state\[8\] vssd1 vssd1 vccd1 vccd1 net1700
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12063__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold176 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 net1711
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 team_01_WB.instance_to_wrap.a1.ADR_I\[18\] vssd1 vssd1 vccd1 vccd1 net1722
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout601 _04754_ vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__buf_2
Xfanout612 net614 vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__buf_4
Xhold198 net105 vssd1 vssd1 vccd1 vccd1 net1733 sky130_fd_sc_hd__dlygate4sd3_1
X_09915_ _06250_ _06253_ vssd1 vssd1 vccd1 vccd1 _06255_ sky130_fd_sc_hd__or2_2
Xfanout623 _04628_ vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__buf_4
XANTENNA__12998__S net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout634 _03733_ vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__clkbuf_2
XANTENNA__14779__A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout675_A _04791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout645 _04839_ vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__clkbuf_2
Xfanout656 _04815_ vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__buf_6
XFILLER_0_42_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11755__X _07941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09846_ _06178_ _06185_ vssd1 vssd1 vccd1 vccd1 _06186_ sky130_fd_sc_hd__or2_2
Xfanout667 _04801_ vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11696__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout678 net679 vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08777__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12893__B1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1003_X net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout689 _04773_ vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_126_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[15\] net812 net773 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[15\]
+ _06116_ vssd1 vssd1 vccd1 vccd1 _06117_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout842_A _03734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13437__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout463_X net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08728_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[5\] net694 _05046_ _05053_
+ _05059_ vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_1_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10656__C1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08659_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[10\] net691 _04986_ _04988_
+ _04991_ vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout630_X net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout728_X net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15403__A net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11670_ net2043 net234 net499 vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__mux2_1
XANTENNA__08943__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10621_ _06886_ _06887_ _06960_ vssd1 vssd1 vccd1 vccd1 _06961_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12238__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08616__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13340_ team_01_WB.instance_to_wrap.cpu.f0.i\[13\] _07679_ net565 vssd1 vssd1 vccd1
+ vccd1 _03815_ sky130_fd_sc_hd__o21ai_1
X_10552_ net505 _06671_ net544 vssd1 vssd1 vccd1 vccd1 _06892_ sky130_fd_sc_hd__mux2_1
XANTENNA__10423__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13271_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[30\] _03761_ net825 vssd1 vssd1
+ vccd1 vccd1 _01898_ sky130_fd_sc_hd__mux2_1
X_10483_ _06781_ _06815_ _06822_ _06818_ vssd1 vssd1 vccd1 vccd1 _06823_ sky130_fd_sc_hd__o31a_1
Xclkbuf_leaf_129_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_129_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15010_ net1350 vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__inv_2
X_12222_ net2066 net290 net444 vssd1 vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__mux2_1
XANTENNA__09577__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13373__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_60_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input69_A wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12153_ net1812 net307 net454 vssd1 vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11104_ _07064_ net327 _07395_ _07443_ vssd1 vssd1 vccd1 vccd1 _07444_ sky130_fd_sc_hd__a22oi_1
XANTENNA__09329__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16961_ clknet_leaf_52_wb_clk_i _02648_ _00944_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_12084_ net1886 net298 net462 vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__mux2_1
XANTENNA__14689__A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13676__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11665__X _07870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11035_ _05006_ _06527_ vssd1 vssd1 vccd1 vccd1 _07375_ sky130_fd_sc_hd__nand2_1
X_15912_ net1399 vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__inv_2
XANTENNA__12701__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16892_ clknet_leaf_59_wb_clk_i _02579_ _00875_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_15843_ net1325 vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__inv_2
X_15774_ net1198 vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__inv_2
X_12986_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[100\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[108\]
+ net860 vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17513_ clknet_leaf_40_wb_clk_i _03200_ _01496_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14725_ net1210 vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__inv_2
XANTENNA__09014__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11937_ net2583 net270 net477 vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__mux2_1
XANTENNA__12937__A _04968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17444_ clknet_leaf_83_wb_clk_i _03131_ _01427_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14656_ net1221 vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__inv_2
X_11868_ net1786 net203 net483 vssd1 vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__mux2_1
XANTENNA__09949__C net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08853__C net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10819_ net530 _07158_ vssd1 vssd1 vccd1 vccd1 _07159_ sky130_fd_sc_hd__nor2_1
X_13607_ net186 _04047_ _04048_ net725 vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__a211o_1
XANTENNA__12939__B2 _03702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17375_ clknet_leaf_44_wb_clk_i _03062_ _01358_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12148__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14587_ net1417 vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__inv_2
X_11799_ net3057 net272 net493 vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__mux2_1
X_16326_ clknet_leaf_93_wb_clk_i _02080_ _00309_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13538_ _03931_ _03990_ vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12943__Y _03705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11987__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13469_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] _05592_ vssd1 vssd1
+ vccd1 vccd1 _03930_ sky130_fd_sc_hd__nand2_1
X_16257_ clknet_leaf_151_wb_clk_i net1627 _00245_ vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15208_ net1382 vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16188_ clknet_leaf_1_wb_clk_i _01948_ _00176_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_58_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15139_ net1220 vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09700_ net1154 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[21\] net953
+ vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__and3_1
XANTENNA__12611__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08543__A1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09631_ net1136 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[23\] net958
+ vssd1 vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_143_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_143_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09562_ _05898_ _05900_ vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14092__A2 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08513_ net1081 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[18\] net940
+ vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_121_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09493_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[30\] net701 _05828_ _05832_
+ vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__o22ai_4
XANTENNA_fanout256_A _07892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08444_ net1004 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[23\] net911
+ vssd1 vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__and3_1
XFILLER_0_65_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08375_ _04626_ _04711_ _04712_ _04714_ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__or4_2
XANTENNA_fanout423_A net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1165_A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13949__Y _04241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09271__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11897__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1332_A net1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17903__1438 vssd1 vssd1 vccd1 vccd1 _17903__1438/HI net1438 sky130_fd_sc_hd__conb_1
XANTENNA__09023__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout792_A net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09891__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1407 net1408 vssd1 vssd1 vccd1 vccd1 net1407 sky130_fd_sc_hd__buf_4
Xfanout420 net422 vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__buf_4
Xfanout1418 net1428 vssd1 vssd1 vccd1 vccd1 net1418 sky130_fd_sc_hd__buf_2
XANTENNA_fanout678_X net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout431 _07964_ vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__buf_6
Xfanout1429 net1430 vssd1 vssd1 vccd1 vccd1 net1429 sky130_fd_sc_hd__clkbuf_4
Xfanout442 _07962_ vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__buf_4
XANTENNA__12521__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout453 _07957_ vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__buf_6
Xfanout464 _07954_ vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout475 _07950_ vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__clkbuf_8
Xfanout486 _07948_ vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__buf_4
XANTENNA__08938__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09829_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[13\] net817 net811 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06169_ sky130_fd_sc_hd__a22o_1
Xfanout497 net498 vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__buf_4
XANTENNA_fanout845_X net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12840_ net2539 net209 net380 vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__mux2_1
XANTENNA__14083__A2 _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12771_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] net1060 net363 _03608_
+ vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__a22o_1
XANTENNA__13860__B net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12094__A1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08837__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11722_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] _07798_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\]
+ vssd1 vssd1 vccd1 vccd1 _07915_ sky130_fd_sc_hd__a21oi_1
X_14510_ net1354 vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15490_ net1321 vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__inv_2
XANTENNA__08673__C net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09131__A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11653_ net719 _07621_ net616 _07859_ vssd1 vssd1 vccd1 vccd1 _07860_ sky130_fd_sc_hd__o211a_1
X_14441_ net1228 vssd1 vssd1 vccd1 vccd1 _00235_ sky130_fd_sc_hd__inv_2
XANTENNA__10277__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09247__C1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09798__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13594__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10604_ _06941_ _06943_ net539 vssd1 vssd1 vccd1 vccd1 _06944_ sky130_fd_sc_hd__mux2_1
X_17160_ clknet_leaf_62_wb_clk_i _02847_ _01143_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_14372_ net1195 vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11584_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] _07800_ vssd1 vssd1 vccd1
+ vccd1 _07801_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09262__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16111_ clknet_leaf_137_wb_clk_i _01886_ _00099_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[18\]
+ sky130_fd_sc_hd__dfrtp_4
X_13323_ _04477_ _03801_ _04518_ vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10535_ _06871_ _06872_ _06873_ _06874_ vssd1 vssd1 vccd1 vccd1 _06875_ sky130_fd_sc_hd__or4_1
X_17091_ clknet_leaf_26_wb_clk_i _02778_ _01074_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13346__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16042_ clknet_leaf_88_wb_clk_i _01836_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13254_ team_01_WB.instance_to_wrap.cpu.f0.i\[23\] _03744_ vssd1 vssd1 vccd1 vccd1
+ _03746_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10466_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[26\] net778 net746 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06806_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12205_ net1839 net267 net443 vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13185_ net25 net837 net630 net2427 vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10397_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[16\] net767 _06730_ _06736_
+ vssd1 vssd1 vccd1 vccd1 _06737_ sky130_fd_sc_hd__o22a_2
Xclkbuf_3_6_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10443__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09970__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12136_ net2252 net270 net451 vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17993_ net1505 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__buf_2
XANTENNA__09009__C net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13649__A2 _07507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12431__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16944_ clknet_leaf_109_wb_clk_i _02631_ _00927_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_12067_ net2033 net204 net459 vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_97_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11018_ _04883_ _06671_ vssd1 vssd1 vccd1 vccd1 _07358_ sky130_fd_sc_hd__xor2_1
XANTENNA__09722__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16875_ clknet_leaf_7_wb_clk_i _02562_ _00858_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_26_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15826_ net1331 vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14074__A2 _04230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13770__B _04146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13282__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15757_ net1341 vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__inv_2
X_12969_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[117\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[125\]
+ net859 vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14708_ net1197 vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15688_ net1376 vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08583__C net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17427_ clknet_leaf_17_wb_clk_i _03114_ _01410_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_14639_ net1291 vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10187__A _06526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09789__A0 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08160_ net1649 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[113\] net1056 vssd1 vssd1
+ vccd1 vccd1 _03527_ sky130_fd_sc_hd__mux2_1
X_17358_ clknet_leaf_28_wb_clk_i _03045_ _01341_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_99_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16309_ clknet_leaf_123_wb_clk_i _02063_ _00292_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08091_ _04525_ _04561_ _04562_ net569 net1541 vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__a32o_1
X_17289_ clknet_leaf_40_wb_clk_i _02976_ _01272_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12606__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload30 clknet_leaf_150_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload30/Y sky130_fd_sc_hd__inv_6
XFILLER_0_24_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload41 clknet_leaf_146_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload41/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_77_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload52 clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload52/Y sky130_fd_sc_hd__bufinv_16
Xclkload63 clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload63/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__10634__B _05835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload74 clknet_leaf_57_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload74/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_51_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload85 clknet_leaf_142_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload85/Y sky130_fd_sc_hd__inv_12
XFILLER_0_11_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload96 clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload96/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_114_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08879__X _05219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10020__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09961__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08993_ net1007 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[8\] net917 vssd1
+ vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_145_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11168__D _07507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12341__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09713__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08758__C net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout373_A _06188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16110__Q team_01_WB.instance_to_wrap.cpu.f0.data_adr\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09614_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[24\] net816 net788 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _05954_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10874__A2 _06811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14065__A2 _04259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09545_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[28\] net783 net753 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[28\]
+ _05871_ vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout638_A _03572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09476_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[30\] net670 net667 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[30\]
+ _05810_ vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10809__B net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08427_ net1116 net1122 net1126 net1120 vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_19_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1070_X net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout805_A net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout426_X net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1168_X net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09886__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08358_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[30\] net821 _04647_ _04679_
+ _04683_ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08790__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload2 clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload2/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12516__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08289_ net1159 net1161 net1164 net1167 vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_150_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13328__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_61_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10320_ net1129 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[18\] net968
+ vssd1 vssd1 vccd1 vccd1 _06660_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout795_X net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10251_ net339 vssd1 vssd1 vccd1 vccd1 _06591_ sky130_fd_sc_hd__inv_2
XANTENNA__10011__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10182_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[10\] net823 net783 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06522_ sky130_fd_sc_hd__a22o_1
XANTENNA__13855__B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1204 net1205 vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__buf_4
Xfanout1215 net1216 vssd1 vssd1 vccd1 vccd1 net1215 sky130_fd_sc_hd__buf_4
Xfanout1226 net1229 vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__buf_4
XANTENNA__12251__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1237 net1242 vssd1 vssd1 vccd1 vccd1 net1237 sky130_fd_sc_hd__clkbuf_4
X_14990_ net1299 vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__inv_2
Xfanout250 _07904_ vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1248 net1303 vssd1 vssd1 vccd1 vccd1 net1248 sky130_fd_sc_hd__buf_2
XANTENNA__08507__A1 net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1259 net1260 vssd1 vssd1 vccd1 vccd1 net1259 sky130_fd_sc_hd__buf_4
Xfanout261 _07880_ vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__buf_2
XANTENNA__08668__C net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09126__A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout272 net275 vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__buf_2
Xfanout283 _07908_ vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__clkbuf_2
X_13941_ _04218_ _04232_ vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__nor2_4
Xfanout294 net295 vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__buf_2
X_16660_ clknet_leaf_67_wb_clk_i _02347_ _00643_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_13872_ net160 net71 net73 vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__and3b_1
XFILLER_0_88_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08965__A net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15611_ net1253 vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__inv_2
X_12823_ net1038 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[3\] vssd1 vssd1 vccd1
+ vccd1 _03645_ sky130_fd_sc_hd__or2_1
X_16591_ clknet_leaf_30_wb_clk_i _02278_ _00574_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[23\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_97_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_141_Right_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15542_ net1261 vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__inv_2
X_12754_ net1034 _07600_ vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__nand2_1
XANTENNA__09483__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11705_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[10\] net714 vssd1 vssd1 vccd1
+ vccd1 _07901_ sky130_fd_sc_hd__or2_1
X_15473_ net1420 vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__inv_2
X_12685_ net3053 net314 net389 vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_144_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_144_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_17212_ clknet_leaf_60_wb_clk_i _02899_ _01195_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11636_ net615 _07846_ _07843_ _07844_ vssd1 vssd1 vccd1 vccd1 _07847_ sky130_fd_sc_hd__a2bb2o_2
X_14424_ net1325 vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09235__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17143_ clknet_leaf_13_wb_clk_i _02830_ _01126_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_14355_ net1333 vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__inv_2
X_11567_ net3095 net154 team_01_WB.instance_to_wrap.cpu.K0.next_state vssd1 vssd1
+ vccd1 vccd1 _03273_ sky130_fd_sc_hd__mux2_1
XANTENNA__10294__X _06634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12426__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10250__A0 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_17 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13319__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10518_ net503 vssd1 vssd1 vccd1 vccd1 _06858_ sky130_fd_sc_hd__inv_2
X_13306_ net566 _07711_ _03788_ net828 vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__a31o_1
XANTENNA__12790__A2 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold709 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[9\] vssd1 vssd1 vccd1 vccd1 net2244
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14286_ net1337 vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__inv_2
X_17074_ clknet_leaf_110_wb_clk_i _02761_ _01057_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11498_ net1683 net876 _07758_ _07776_ vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_94_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16025_ net1324 vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__inv_2
X_13237_ net2636 net354 net350 team_01_WB.instance_to_wrap.cpu.f0.i\[13\] vssd1 vssd1
+ vccd1 vccd1 _01913_ sky130_fd_sc_hd__a22o_1
X_10449_ net1147 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[26\] net979
+ vssd1 vssd1 vccd1 vccd1 _06789_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13168_ net2363 net848 net840 net1974 vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12119_ net2862 net311 net458 vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__mux2_1
XANTENNA__12161__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13099_ _03719_ _03720_ _03721_ _03722_ vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__or4_1
X_17976_ net1491 vssd1 vssd1 vccd1 vccd1 la_data_out[18] sky130_fd_sc_hd__buf_2
Xhold1409 _03512_ vssd1 vssd1 vccd1 vccd1 net2944 sky130_fd_sc_hd__dlygate4sd3_1
X_16927_ clknet_leaf_43_wb_clk_i _02614_ _00910_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11285__B _07566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16858_ clknet_leaf_76_wb_clk_i _02545_ _00841_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14047__A2 _04226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17902__1437 vssd1 vssd1 vccd1 vccd1 _17902__1437/HI net1437 sky130_fd_sc_hd__conb_1
X_15809_ net1197 vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_49_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16789_ clknet_leaf_114_wb_clk_i _02476_ _00772_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10469__X _06809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09330_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[24\] net675 net667 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_46_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09261_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[20\] net692 net674 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_66_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09202__C net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10348__C net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08212_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[69\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[61\]
+ net1050 vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09192_ net1087 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[17\] net923
+ vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09226__A2 _05564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08143_ _04479_ team_01_WB.instance_to_wrap.cpu.f0.num\[15\] _04498_ team_01_WB.instance_to_wrap.cpu.f0.i\[2\]
+ _04589_ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_116_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12336__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout219_A net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10241__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload130 clknet_leaf_79_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload130/Y sky130_fd_sc_hd__inv_6
XANTENNA__12781__A2 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08074_ _04524_ _04547_ vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__nand2_1
Xclkload141 clknet_leaf_81_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload141/Y sky130_fd_sc_hd__inv_12
XANTENNA__10792__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08115__A team_01_WB.instance_to_wrap.cpu.f0.i\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16105__Q team_01_WB.instance_to_wrap.cpu.f0.data_adr\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1030_A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1128_A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09934__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13730__B2 net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout490_A _07947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12071__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 net145 vssd1 vssd1 vccd1 vccd1 net1549 sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ net1087 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[8\] net917 vssd1
+ vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__and3_1
Xhold25 _02023_ vssd1 vssd1 vccd1 vccd1 net1560 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09147__D1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold36 team_01_WB.instance_to_wrap.cpu.f0.write_data\[5\] vssd1 vssd1 vccd1 vccd1
+ net1571 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13962__Y _04254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold47 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[4\] vssd1 vssd1 vccd1 vccd1 net1582
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net1593 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_85_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold69 net88 vssd1 vssd1 vccd1 vccd1 net1604 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout755_A _04675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout376_X net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08785__A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout922_A _04770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09528_ _05805_ _05807_ vssd1 vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09465__A2 _05803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09459_ _05784_ _05796_ _05797_ _05798_ vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout808_X net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13549__A1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12470_ net2335 net234 net411 vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__mux2_1
XANTENNA__09217__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12754__B _07600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11421_ net323 _07733_ _07734_ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__and3_1
XFILLER_0_152_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12246__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10555__A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10232__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14140_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[95\] _04241_ _04256_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[47\]
+ vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11352_ _04481_ _07680_ vssd1 vssd1 vccd1 vccd1 _07681_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10303_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[18\] net754 net752 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06643_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14071_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[68\] _04247_ _04253_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__a22o_1
X_11283_ _07188_ _07232_ _07553_ _07600_ vssd1 vssd1 vccd1 vccd1 _07623_ sky130_fd_sc_hd__or4b_1
XFILLER_0_46_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13022_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[64\] net2801 net857 vssd1 vssd1
+ vccd1 vccd1 _02103_ sky130_fd_sc_hd__mux2_1
X_10234_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[9\] net797 net791 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06574_ sky130_fd_sc_hd__a22o_1
XANTENNA_input51_A wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11732__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1001 net1002 vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__clkbuf_2
Xfanout1012 net1013 vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11386__A team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17830_ clknet_leaf_119_wb_clk_i _03506_ _01770_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[100\]
+ sky130_fd_sc_hd__dfstp_1
X_10165_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[10\] net803 net732 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[10\]
+ _06504_ vssd1 vssd1 vccd1 vccd1 _06505_ sky130_fd_sc_hd__a221o_1
XANTENNA__10290__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1023 net1024 vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__buf_1
Xfanout1034 team_01_WB.instance_to_wrap.cpu.RU0.InstrRead vssd1 vssd1 vccd1 vccd1
+ net1034 sky130_fd_sc_hd__clkbuf_4
Xfanout1045 net1059 vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__clkbuf_4
Xfanout1056 net1058 vssd1 vssd1 vccd1 vccd1 net1056 sky130_fd_sc_hd__clkbuf_4
X_17761_ clknet_leaf_121_wb_clk_i _03437_ _01701_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10096_ _06426_ _06430_ _06435_ vssd1 vssd1 vccd1 vccd1 _06436_ sky130_fd_sc_hd__or3_4
Xfanout1067 team_01_WB.instance_to_wrap.cpu.RU0.state\[4\] vssd1 vssd1 vccd1 vccd1
+ net1067 sky130_fd_sc_hd__buf_2
X_14973_ net1311 vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__inv_2
Xfanout1078 net1079 vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__buf_1
XFILLER_0_156_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1089 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[24\] vssd1 vssd1 vccd1 vccd1
+ net1089 sky130_fd_sc_hd__clkbuf_2
X_16712_ clknet_leaf_27_wb_clk_i _02399_ _00695_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13924_ net2906 _04215_ _04216_ vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__o21a_1
XANTENNA__10838__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17692_ clknet_leaf_137_wb_clk_i _03376_ _01633_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__14029__A2 _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12929__B net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16643_ clknet_leaf_28_wb_clk_i _02330_ _00626_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13855_ net1180 net1067 net1655 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[16\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_53_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13106__A net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12806_ net1998 net640 net608 _03632_ vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__a22o_1
X_16574_ clknet_leaf_115_wb_clk_i _02261_ _00557_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_13786_ _04158_ _04169_ vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__nand2_1
X_10998_ net558 _05263_ _06902_ vssd1 vssd1 vccd1 vccd1 _07338_ sky130_fd_sc_hd__or3_1
XANTENNA__09456__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15525_ net1288 vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09022__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12737_ net1862 net638 net606 _03585_ vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_26_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10471__B1 _06809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15456_ net1234 vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12668_ net2231 net233 net387 vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09957__C net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08861__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14407_ net1358 vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__inv_2
XANTENNA__12156__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11619_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] _07819_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\]
+ vssd1 vssd1 vccd1 vccd1 _07833_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_61_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15387_ net1253 vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__inv_2
X_12599_ net3109 net242 net397 vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_133_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17126_ clknet_leaf_73_wb_clk_i _02813_ _01109_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14338_ net1338 vssd1 vssd1 vccd1 vccd1 _00132_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold506 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2041 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10184__B net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold517 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[21\] vssd1 vssd1 vccd1 vccd1
+ net2052 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11995__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold528 team_01_WB.instance_to_wrap.cpu.f0.write_data\[7\] vssd1 vssd1 vccd1 vccd1
+ net2063 sky130_fd_sc_hd__dlygate4sd3_1
X_17057_ clknet_leaf_55_wb_clk_i _02744_ _01040_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold539 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2074 sky130_fd_sc_hd__dlygate4sd3_1
X_14269_ net1204 vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__inv_2
XANTENNA__09916__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16008_ net1357 vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_41_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11296__A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08830_ net1104 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[1\] net938 vssd1
+ vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__and3_1
XFILLER_0_148_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1206 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2741 sky130_fd_sc_hd__dlygate4sd3_1
X_08761_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[4\] net656 _05084_ _05095_
+ _05098_ vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__a2111o_1
Xhold1217 team_01_WB.instance_to_wrap.cpu.f0.num\[21\] vssd1 vssd1 vccd1 vccd1 net2752
+ sky130_fd_sc_hd__dlygate4sd3_1
X_17959_ net1474 vssd1 vssd1 vccd1 vccd1 la_data_out[1] sky130_fd_sc_hd__buf_2
Xhold1228 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2763 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1239 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[47\] vssd1 vssd1 vccd1 vccd1
+ net2774 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08692_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[7\] net680 _05009_ _05011_
+ _05016_ vssd1 vssd1 vccd1 vccd1 _05032_ sky130_fd_sc_hd__a2111o_1
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_105_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09447__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09313_ _05649_ _05650_ _05651_ _05652_ vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_24_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout336_A net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10078__C net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1078_A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10462__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09244_ _05572_ _05581_ _05582_ _05583_ vssd1 vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__or4_1
XANTENNA_wire978_X net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08771__C net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09175_ net1010 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[16\] net944
+ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13400__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12066__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout503_A _06857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1245_A net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08126_ _04473_ team_01_WB.instance_to_wrap.cpu.f0.num\[21\] team_01_WB.instance_to_wrap.cpu.f0.num\[17\]
+ _04477_ vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13957__Y _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10765__A1 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08057_ team_01_WB.instance_to_wrap.cpu.f0.i\[6\] team_01_WB.instance_to_wrap.cpu.K0.keyvalid
+ _04523_ _04534_ vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout1033_X net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout872_A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout493_X net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13973__X _04265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1200_X net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11190__A1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08959_ _05290_ _05291_ _05297_ _05298_ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout660_X net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout758_X net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12809__A3 _03634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11970_ net2170 net243 net473 vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__mux2_1
XANTENNA__09686__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08946__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10921_ net522 _07218_ _07150_ _07040_ vssd1 vssd1 vccd1 vccd1 _07261_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout925_X net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10852_ _06501_ _06530_ _07191_ vssd1 vssd1 vccd1 vccd1 _07192_ sky130_fd_sc_hd__or3_1
X_13640_ net987 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] _04075_ _04076_
+ vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12442__A1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13571_ net986 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] _04017_ _04018_
+ vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__a22o_1
X_10783_ _06944_ _06950_ net520 vssd1 vssd1 vccd1 vccd1 _07123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15310_ net1291 vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__inv_2
X_12522_ _07793_ _07951_ net573 vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__and3_1
X_16290_ clknet_leaf_100_wb_clk_i _02044_ _00273_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[13\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_136_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08681__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15241_ net1288 vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__inv_2
X_12453_ net2311 net317 net418 vssd1 vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12745__A2 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11404_ _07695_ net323 _07725_ vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__and3b_1
X_12384_ net2024 net292 net426 vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15172_ net1230 vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09610__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11335_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[1\] net1176 _04559_ _07652_ vssd1
+ vssd1 vccd1 vccd1 _07666_ sky130_fd_sc_hd__a22o_1
X_14123_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[14\] _04253_ _04256_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[46\]
+ vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__a22o_1
XANTENNA__10572__X _06912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17901__1436 vssd1 vssd1 vccd1 vccd1 _17901__1436/HI net1436 sky130_fd_sc_hd__conb_1
XANTENNA__12704__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11266_ net374 net333 net331 vssd1 vssd1 vccd1 vccd1 _07606_ sky130_fd_sc_hd__a21o_1
X_14054_ _04236_ _04247_ _04258_ _04259_ vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__or4_1
XANTENNA__10732__B _05898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10217_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[8\] net793 net736 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _06557_ sky130_fd_sc_hd__a22o_1
X_13005_ net3000 net2935 net866 vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11197_ _05529_ net331 _07536_ net369 vssd1 vssd1 vccd1 vccd1 _07537_ sky130_fd_sc_hd__a211o_1
XFILLER_0_101_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10451__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17813_ clknet_leaf_95_wb_clk_i net2408 _01753_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[83\]
+ sky130_fd_sc_hd__dfrtp_1
X_10148_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[11\] net801 net755 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06488_ sky130_fd_sc_hd__a22o_1
XANTENNA__09017__C net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17744_ clknet_leaf_116_wb_clk_i _03420_ _01684_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14956_ net1260 vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__inv_2
X_10079_ net1138 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[7\] net954 vssd1
+ vssd1 vccd1 vccd1 _06419_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09677__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13907_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[7\] _04204_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__a21o_1
X_17675_ clknet_leaf_0_wb_clk_i _03360_ _01616_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_14887_ net1390 vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__inv_2
X_16626_ clknet_leaf_143_wb_clk_i _02313_ _00609_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13838_ net1615 net830 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[31\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_98_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09429__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12946__Y _03707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12433__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16557_ clknet_leaf_157_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[23\]
+ _00540_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13769_ _04156_ vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_63_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15051__A net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15508_ net1380 vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__inv_2
X_16488_ clknet_leaf_152_wb_clk_i _02242_ _00471_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10995__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15439_ net1386 vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_152_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12736__A2 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold303 team_01_WB.instance_to_wrap.a1.ADR_I\[26\] vssd1 vssd1 vccd1 vccd1 net1838
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold314 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[31\] vssd1 vssd1 vccd1 vccd1 net1849
+ sky130_fd_sc_hd__dlygate4sd3_1
X_17109_ clknet_leaf_110_wb_clk_i _02796_ _01092_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold325 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1860 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12614__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold336 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1871 sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net1882 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold358 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1893 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[4\] net780 net748 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06271_ sky130_fd_sc_hd__a22o_1
Xhold369 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[21\] vssd1 vssd1 vccd1 vccd1 net1904
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout805 net806 vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_21_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout816 _04636_ vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09365__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13161__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09862_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[12\] net816 net770 _06196_
+ vssd1 vssd1 vccd1 vccd1 _06202_ sky130_fd_sc_hd__a211o_1
Xfanout827 _04579_ vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__clkbuf_4
Xfanout838 _03736_ vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__buf_1
Xfanout849 net850 vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__clkbuf_2
X_08813_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\] net729 vssd1 vssd1 vccd1 vccd1
+ _05153_ sky130_fd_sc_hd__and2_1
Xhold1003 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[59\] vssd1 vssd1 vccd1 vccd1
+ net2538 sky130_fd_sc_hd__dlygate4sd3_1
X_09793_ net374 _06131_ vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__nor2_1
Xhold1014 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1025 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2560 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout286_A _07896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1036 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1047 team_01_WB.instance_to_wrap.cpu.f0.num\[12\] vssd1 vssd1 vccd1 vccd1 net2582
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08744_ net1099 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[4\] net880 vssd1
+ vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__and3_1
Xhold1058 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2593 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_107_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1069 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2604 sky130_fd_sc_hd__dlygate4sd3_1
X_08675_ net1085 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[7\] net926 vssd1
+ vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout453_A _07957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09878__B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1362_A net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout718_A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout339_X net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09597__C net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09840__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09227_ _05529_ _05566_ vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_8_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1248_X net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09158_ net1017 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[16\] net904
+ vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08109_ _04504_ net1176 vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__nand2_2
X_09089_ net1094 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[13\] net918
+ vssd1 vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12524__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11120_ _06313_ net334 net332 vssd1 vssd1 vccd1 vccd1 _07460_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold870 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold881 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2416 sky130_fd_sc_hd__dlygate4sd3_1
Xhold892 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 net2427
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13152__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11051_ _07389_ _07390_ _07388_ vssd1 vssd1 vccd1 vccd1 _07391_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08022__B _04516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10002_ net516 _06341_ vssd1 vssd1 vccd1 vccd1 _06342_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10271__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14810_ net1371 vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15790_ net1190 vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__inv_2
XANTENNA__08676__C net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1570 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net3105 sky130_fd_sc_hd__dlygate4sd3_1
X_14741_ net1194 vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__inv_2
XANTENNA_input14_A DAT_I[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1581 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1592 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net3127 sky130_fd_sc_hd__dlygate4sd3_1
X_11953_ net2563 net311 net477 vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10904_ net335 _07243_ vssd1 vssd1 vccd1 vccd1 _07244_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_84_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17460_ clknet_leaf_22_wb_clk_i _03147_ _01443_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_14672_ net1307 vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__inv_2
X_11884_ net2652 net278 net483 vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16411_ clknet_leaf_125_wb_clk_i _02165_ _00394_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13623_ net989 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] _04061_ _04062_
+ vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11218__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10835_ _06193_ _06218_ _07173_ _06192_ _06164_ vssd1 vssd1 vccd1 vccd1 _07175_ sky130_fd_sc_hd__a311oi_4
XANTENNA__08619__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17391_ clknet_leaf_34_wb_clk_i _03078_ _01374_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13090__S net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16342_ clknet_leaf_93_wb_clk_i net2598 _00325_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[65\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13554_ net720 _07621_ net1073 vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__o21a_1
X_10766_ _07104_ _07105_ net520 vssd1 vssd1 vccd1 vccd1 _07106_ sky130_fd_sc_hd__mux2_1
XANTENNA__09831__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10977__A1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12505_ net2102 net263 net407 vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__mux2_1
X_16273_ clknet_leaf_88_wb_clk_i _00001_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA__09300__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13485_ _03850_ _03851_ _03943_ _03848_ _03847_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__a311o_1
X_10697_ _06941_ _06949_ net535 vssd1 vssd1 vccd1 vccd1 _07037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18012_ net637 vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10446__C net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15224_ net1212 vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__inv_2
X_12436_ net3162 net238 net415 vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15155_ net1405 vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12367_ net1970 net200 net423 vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12434__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14215__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[17\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14106_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[37\] _04230_ _04255_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[117\]
+ _04392_ vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__a221o_1
X_11318_ _04505_ _07652_ _07654_ _07650_ vssd1 vssd1 vccd1 vccd1 _07655_ sky130_fd_sc_hd__a211o_4
X_15086_ net1298 vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12298_ net3121 net207 net433 vssd1 vssd1 vccd1 vccd1 _02696_ sky130_fd_sc_hd__mux2_1
XANTENNA__13143__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14037_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[2\] _04265_ _04289_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[2\]
+ _04152_ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__a221o_1
X_11249_ _07588_ vssd1 vssd1 vccd1 vccd1 _07589_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_56_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09898__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_max_cap304_X net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15988_ net1368 vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__inv_2
XANTENNA__08586__C net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17727_ clknet_leaf_150_wb_clk_i _03404_ _01668_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_14939_ net1274 vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08460_ net1025 net889 vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__and2_2
X_17658_ clknet_leaf_3_wb_clk_i net1667 _01599_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_102_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16609_ clknet_leaf_50_wb_clk_i _02296_ _00592_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_08391_ _04724_ _04730_ vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__nand2_1
X_17589_ clknet_leaf_130_wb_clk_i _03276_ _01548_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.code\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12609__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11513__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09210__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09012_ net1099 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[9\] net943 vssd1
+ vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold100 _02009_ vssd1 vssd1 vccd1 vccd1 net1635 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12344__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold111 team_01_WB.instance_to_wrap.cpu.f0.write_data\[18\] vssd1 vssd1 vccd1 vccd1
+ net1646 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout201_A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold122 _01970_ vssd1 vssd1 vccd1 vccd1 net1657 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_84 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold133 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 net1668
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 _01993_ vssd1 vssd1 vccd1 vccd1 net1679 sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 _01973_ vssd1 vssd1 vccd1 vccd1 net1690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 net1701
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold177 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[20\] vssd1 vssd1 vccd1 vccd1
+ net1712 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16113__Q team_01_WB.instance_to_wrap.cpu.f0.data_adr\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold188 _02016_ vssd1 vssd1 vccd1 vccd1 net1723 sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 _02006_ vssd1 vssd1 vccd1 vccd1 net1734 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13134__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout602 net603 vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__buf_4
X_09914_ _06250_ _06253_ vssd1 vssd1 vccd1 vccd1 _06254_ sky130_fd_sc_hd__nand2_1
Xfanout613 net614 vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1110_A net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout624 _04628_ vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout635 net636 vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1208_A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout646 _04825_ vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__clkbuf_8
X_09845_ _06180_ _06182_ _06183_ _06184_ vssd1 vssd1 vccd1 vccd1 _06185_ sky130_fd_sc_hd__or4_1
Xfanout657 _04815_ vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__buf_4
XANTENNA_input6_A DAT_I[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout668 _04801_ vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__buf_4
XANTENNA__12893__A1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11696__A2 _07520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout679 _04789_ vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__buf_8
XANTENNA_fanout668_A _04801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14095__B1 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09776_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[15\] net805 net746 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06116_ sky130_fd_sc_hd__a22o_1
XANTENNA__13970__Y _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08727_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[5\] net692 _05054_ _05056_
+ _05062_ vssd1 vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12867__X _03652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08849__B1 _05188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout456_X net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout835_A _03737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09889__A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08658_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[10\] net697 _04978_
+ _04979_ _04990_ vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10120__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17900__1435 vssd1 vssd1 vccd1 vccd1 _17900__1435/HI net1435 sky130_fd_sc_hd__conb_1
XFILLER_0_96_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout623_X net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12519__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08589_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[15\] net691 net658 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10620_ _06934_ _06959_ _06927_ _06933_ vssd1 vssd1 vccd1 vccd1 _06960_ sky130_fd_sc_hd__a211o_1
XANTENNA__12948__A2 _03707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10551_ _06707_ net371 net544 vssd1 vssd1 vccd1 vccd1 _06891_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09120__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10266__C net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13858__B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13270_ net587 _03750_ _03759_ _03760_ vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__a31o_1
X_10482_ _06814_ _06820_ vssd1 vssd1 vccd1 vccd1 _06822_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11659__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12221_ net2487 net313 net445 vssd1 vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__mux2_1
XANTENNA__12254__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12152_ net2272 net311 net452 vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__mux2_1
XANTENNA__09129__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11103_ net556 _06280_ net334 _07442_ vssd1 vssd1 vccd1 vccd1 _07443_ sky130_fd_sc_hd__a31o_1
XANTENNA__13125__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16960_ clknet_leaf_46_wb_clk_i _02647_ _00943_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_12083_ net1877 net276 net459 vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11034_ _04969_ net340 vssd1 vssd1 vccd1 vccd1 _07374_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09416__X _05756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15911_ net1412 vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_34_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16891_ clknet_leaf_70_wb_clk_i _02578_ _00874_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12884__A1 _03663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08320__X _04660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15842_ net1326 vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ net1199 vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12985_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[101\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[109\]
+ net859 vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17512_ clknet_leaf_64_wb_clk_i _03199_ _01495_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14724_ net1209 vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11936_ net2366 net241 net477 vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__mux2_1
XANTENNA__10111__A2 _04649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12937__B _07756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17443_ clknet_leaf_29_wb_clk_i _03130_ _01426_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14655_ net1320 vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__inv_2
X_11867_ net2513 net273 net485 vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__mux2_1
XANTENNA__12429__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13606_ net197 net193 _07807_ _07895_ net643 vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__o2111a_1
XPHY_EDGE_ROW_151_Left_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17374_ clknet_leaf_85_wb_clk_i _03061_ _01357_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10818_ _07156_ _07157_ net519 vssd1 vssd1 vccd1 vccd1 _07158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14586_ net1366 vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__inv_2
XANTENNA__09265__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09804__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11798_ net2075 net206 net493 vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16325_ clknet_leaf_120_wb_clk_i net2389 _00308_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13537_ _03925_ _03935_ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10749_ _06744_ _06747_ _06106_ vssd1 vssd1 vccd1 vccd1 _07089_ sky130_fd_sc_hd__a21o_1
XFILLER_0_131_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16256_ clknet_leaf_156_wb_clk_i net1723 _00244_ vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14010__B1 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13468_ _03926_ _03928_ vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__and2_1
XFILLER_0_140_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15207_ net1396 vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__inv_2
X_12419_ net2691 net305 net422 vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16187_ clknet_leaf_1_wb_clk_i _01947_ _00175_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12164__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10178__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13399_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\]
+ net595 vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11288__B team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15138_ net1351 vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__inv_2
XANTENNA__13116__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15069_ net1313 vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_75_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12875__A1 _03657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_155_Right_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08543__A2 _04881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09630_ net1136 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[23\] net951
+ vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_143_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09561_ _05898_ _05900_ vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__nand2_1
XANTENNA__09205__C net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12687__X _03570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08884__Y _05224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08512_ net1001 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[18\] net925 vssd1
+ vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_121_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_121_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09492_ _05816_ _05819_ _05830_ _05831_ vssd1 vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__or4_2
XANTENNA__17699__Q team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_66_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08443_ net1027 net912 vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__and2_1
XANTENNA__12339__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout249_A _07904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08374_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] net1169 vssd1 vssd1 vccd1
+ vccd1 _04714_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16108__Q team_01_WB.instance_to_wrap.cpu.f0.data_adr\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1060_A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout416_A _03562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire960_X net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1158_A net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14001__B1 _04254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13355__A2 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12074__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10169__A2 _04654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout785_A net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1113_X net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11118__A1 _06928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1408 net1409 vssd1 vssd1 vccd1 vccd1 net1408 sky130_fd_sc_hd__clkbuf_4
Xfanout410 _03564_ vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__buf_4
Xfanout1419 net1422 vssd1 vssd1 vccd1 vccd1 net1419 sky130_fd_sc_hd__buf_4
Xfanout421 net422 vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__buf_6
Xfanout432 _07964_ vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13512__C1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout443 _07959_ vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__buf_6
Xfanout454 _07957_ vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12866__A1 net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout952_A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout465 _07954_ vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__buf_6
Xfanout476 _07950_ vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08534__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09828_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[13\] net799 net734 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06168_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout487 _07947_ vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__buf_6
Xfanout498 _07943_ vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__buf_6
XANTENNA_fanout740_X net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09759_ _05618_ _05731_ vssd1 vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09495__A0 _05833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12770_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[19\] _07135_ net1034 vssd1 vssd1
+ vccd1 vccd1 _03608_ sky130_fd_sc_hd__mux2_1
XANTENNA__13291__A1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11721_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[7\] net714 net616 vssd1 vssd1
+ vccd1 vccd1 _07914_ sky130_fd_sc_hd__o21a_1
XANTENNA__12249__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14440_ net1307 vssd1 vssd1 vccd1 vccd1 _00234_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11652_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[21\] net713 vssd1 vssd1 vccd1
+ vccd1 _07859_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10603_ net550 _06496_ _06942_ vssd1 vssd1 vccd1 vccd1 _06943_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13594__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14371_ net1195 vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11583_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\]
+ _07798_ vssd1 vssd1 vccd1 vccd1 _07800_ sky130_fd_sc_hd__and3_1
X_16110_ clknet_leaf_137_wb_clk_i _01885_ _00098_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[17\]
+ sky130_fd_sc_hd__dfrtp_4
X_13322_ net610 _07703_ vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17090_ clknet_leaf_78_wb_clk_i _02777_ _01073_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10534_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[31\] net698 net679 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06874_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16041_ clknet_leaf_88_wb_clk_i _01835_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13253_ _03744_ vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__inv_2
X_10465_ _06801_ _06802_ _06803_ _06804_ vssd1 vssd1 vccd1 vccd1 _06805_ sky130_fd_sc_hd__or4_1
XFILLER_0_150_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12204_ net2299 net234 net443 vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__mux2_1
X_10396_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[16\] net791 _06731_
+ _06734_ _06735_ vssd1 vssd1 vccd1 vccd1 _06736_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_20_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13184_ net26 net835 net628 net1615 vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__o22a_1
XFILLER_0_86_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12135_ net1968 net242 net453 vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__mux2_1
X_17992_ net635 vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12712__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11109__A1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16943_ clknet_leaf_34_wb_clk_i _02630_ _00926_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_12066_ net2905 net273 net461 vssd1 vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__mux2_1
X_11017_ _07355_ _07356_ _07353_ vssd1 vssd1 vccd1 vccd1 _07357_ sky130_fd_sc_hd__and3b_1
X_16874_ clknet_leaf_11_wb_clk_i _02561_ _00857_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_15825_ net1202 vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15324__A net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15756_ net1341 vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12968_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[118\] net1875 net855 vssd1 vssd1
+ vccd1 vccd1 _02157_ sky130_fd_sc_hd__mux2_1
XANTENNA__09486__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_36_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_66_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08864__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14707_ net1193 vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__inv_2
X_11919_ net2303 net294 net481 vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__mux2_1
X_15687_ net1390 vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__inv_2
XANTENNA__12159__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12899_ net356 _03673_ _03674_ net869 net1587 vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__a32o_1
X_17426_ clknet_leaf_144_wb_clk_i _03113_ _01409_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14638_ net1393 vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__inv_2
XANTENNA__09238__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09789__A1 _06128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11998__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17357_ clknet_leaf_67_wb_clk_i _03044_ _01340_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_14569_ net1413 vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12793__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16308_ clknet_leaf_120_wb_clk_i _02062_ _00291_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_08090_ team_01_WB.instance_to_wrap.cpu.f0.i\[0\] _04524_ vssd1 vssd1 vccd1 vccd1
+ _04562_ sky130_fd_sc_hd__or2_1
X_17288_ clknet_leaf_63_wb_clk_i _02975_ _01271_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload20 clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload20/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_77_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16239_ clknet_leaf_141_wb_clk_i net1638 _00227_ vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__dfrtp_1
Xclkload31 clknet_leaf_151_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload31/Y sky130_fd_sc_hd__clkinv_2
Xclkload42 clknet_leaf_147_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload42/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_77_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload53 clknet_leaf_44_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload53/Y sky130_fd_sc_hd__inv_6
XFILLER_0_24_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload64 clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload64/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_149_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload75 clknet_leaf_58_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload75/Y sky130_fd_sc_hd__bufinv_16
Xclkload86 clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload86/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__09410__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload97 clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload97/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_11_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08104__C _04574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12622__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08992_ net1007 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[8\] net882 vssd1
+ vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_145_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10931__A _05338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_75_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10859__A0 _06129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10323__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09613_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[24\] net761 net751 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[24\]
+ _05940_ vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__a221o_1
X_17914__1445 vssd1 vssd1 vccd1 vccd1 _17914__1445/HI net1445 sky130_fd_sc_hd__conb_1
XANTENNA__10874__A3 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09544_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[28\] net809 net751 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__a22o_1
XANTENNA__09477__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12069__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09475_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[30\] net897
+ vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout533_A _05190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_920 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08426_ net1115 net933 vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__and2_2
XFILLER_0_108_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout700_A _04760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08357_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[30\] net815 net794 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload3 clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload3/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA_fanout419_X net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12784__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08288_ _04625_ _04626_ vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__or2_4
XANTENNA__10825__B net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13976__X _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10250_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] _06589_ net623 vssd1
+ vssd1 vccd1 vccd1 _06590_ sky130_fd_sc_hd__mux2_2
XANTENNA_fanout690_X net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09401__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout788_X net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10181_ _06503_ _06519_ _06520_ vssd1 vssd1 vccd1 vccd1 _06521_ sky130_fd_sc_hd__nor3_1
XFILLER_0_121_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12532__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1205 net1206 vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08949__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1216 net1223 vssd1 vssd1 vccd1 vccd1 net1216 sky130_fd_sc_hd__clkbuf_2
Xfanout1227 net1229 vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10560__B _04743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout240 _07870_ vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout955_X net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1238 net1241 vssd1 vssd1 vccd1 vccd1 net1238 sky130_fd_sc_hd__buf_4
Xfanout251 _07904_ vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__clkbuf_2
Xfanout1249 net1252 vssd1 vssd1 vccd1 vccd1 net1249 sky130_fd_sc_hd__buf_4
Xfanout262 _07880_ vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__buf_1
Xfanout273 net275 vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__buf_2
X_13940_ _04228_ _04231_ vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__nand2_2
Xfanout284 _07896_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__buf_2
XANTENNA__11511__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout295 _07926_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__dlymetal6s2s_1
X_13871_ net1536 net1182 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.next_keyvalid
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15610_ net1370 vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__inv_2
X_12822_ net1037 _07464_ vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__nand2_1
XANTENNA__13264__A1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16590_ clknet_leaf_28_wb_clk_i _02277_ _00573_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[22\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_69_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08684__C net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15541_ net1276 vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__inv_2
XANTENNA__11275__B1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12753_ net1559 net640 net608 _03596_ vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14983__A net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11704_ net2267 net226 net499 vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__mux2_1
X_15472_ net1282 vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__inv_2
XANTENNA__08981__A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12684_ net2060 net317 net390 vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17211_ clknet_leaf_70_wb_clk_i _02898_ _01194_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14423_ net1308 vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11635_ _07818_ _07845_ vssd1 vssd1 vccd1 vccd1 _07846_ sky130_fd_sc_hd__or2_1
XANTENNA__12707__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11611__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12775__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17142_ clknet_leaf_30_wb_clk_i _02829_ _01125_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14354_ net1333 vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__inv_2
X_11566_ team_01_WB.instance_to_wrap.cpu.K0.count\[0\] team_01_WB.instance_to_wrap.cpu.K0.count\[1\]
+ vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__nand2b_1
XFILLER_0_64_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13305_ _04473_ _07709_ vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__nand2_1
XANTENNA__10250__A1 _06589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10517_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[31\] net625 _06855_ _06856_
+ vssd1 vssd1 vccd1 vccd1 _06857_ sky130_fd_sc_hd__a22o_2
XANTENNA__13111__B net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17073_ clknet_leaf_116_wb_clk_i _02760_ _01056_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_14285_ net1336 vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11497_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[14\] _07756_ vssd1 vssd1 vccd1
+ vccd1 _07776_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_113_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_113_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10454__C net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16024_ net1324 vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_94_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13236_ net2683 net354 net350 team_01_WB.instance_to_wrap.cpu.f0.i\[14\] vssd1 vssd1
+ vccd1 vccd1 _01914_ sky130_fd_sc_hd__a22o_1
X_10448_ net1147 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[26\] net952
+ vssd1 vssd1 vccd1 vccd1 _06788_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15319__A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12442__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13167_ net1899 net848 net840 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[9\] vssd1
+ vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__a22o_1
X_10379_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[16\] net790 net749 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06719_ sky130_fd_sc_hd__a22o_1
X_12118_ net1750 net294 net458 vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__mux2_1
XANTENNA__08859__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17975_ net1490 vssd1 vssd1 vccd1 vccd1 la_data_out[17] sky130_fd_sc_hd__buf_2
X_13098_ net43 net42 net45 net44 vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__or4_1
X_16926_ clknet_leaf_85_wb_clk_i _02613_ _00909_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12049_ net1853 net301 net464 vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__mux2_1
XANTENNA__10305__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16857_ clknet_leaf_104_wb_clk_i _02544_ _00840_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_159_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11582__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15808_ net1207 vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__inv_2
X_16788_ clknet_leaf_67_wb_clk_i _02475_ _00771_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11266__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15739_ net1254 vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09260_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[20\] net688 net678 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_66_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08211_ net2723 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[62\] net1043 vssd1 vssd1
+ vccd1 vccd1 _03476_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_138_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17409_ clknet_leaf_60_wb_clk_i _03096_ _01392_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_09191_ net1004 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[17\] net939 vssd1
+ vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__and3_1
XANTENNA__12617__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08142_ _04474_ team_01_WB.instance_to_wrap.cpu.f0.num\[20\] team_01_WB.instance_to_wrap.cpu.f0.num\[7\]
+ _04486_ _04597_ vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_116_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08073_ _04525_ _04548_ _04549_ net570 net1571 vssd1 vssd1 vccd1 vccd1 _03541_ sky130_fd_sc_hd__a32o_1
Xclkload120 clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload120/Y sky130_fd_sc_hd__inv_8
Xclkload131 clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload131/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_102_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload142 clknet_leaf_83_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload142/Y sky130_fd_sc_hd__inv_8
XFILLER_0_114_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_842 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13191__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12352__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1023_A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08975_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[8\] net674 _05312_ _05313_
+ _05314_ vssd1 vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__a2111oi_1
Xhold15 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[0\] vssd1 vssd1 vccd1 vccd1
+ net1550 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout483_A _07948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold26 net159 vssd1 vssd1 vccd1 vccd1 net1561 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[5\] vssd1 vssd1 vccd1 vccd1
+ net1572 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16121__Q team_01_WB.instance_to_wrap.cpu.f0.data_adr\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold48 team_01_WB.instance_to_wrap.cpu.LCD0.lcd_rs vssd1 vssd1 vccd1 vccd1 net1583
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 net116 vssd1 vssd1 vccd1 vccd1 net1594 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout650_A _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout369_X net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13246__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09527_ net583 _05866_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] net627
+ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout1180_X net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout915_A net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09458_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[29\] _04766_ net677
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[29\] vssd1 vssd1 vccd1 vccd1
+ _05798_ sky130_fd_sc_hd__a22o_1
XANTENNA__09870__B1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_958 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08409_ _04738_ _04745_ _04736_ vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__and3b_1
XFILLER_0_149_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout703_X net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09389_ net598 _05726_ _05728_ vssd1 vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__o21ai_2
XANTENNA__12527__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11420_ team_01_WB.instance_to_wrap.cpu.f0.i\[16\] _07704_ _07700_ vssd1 vssd1 vccd1
+ vccd1 _07734_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_980 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09622__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08306__A net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10555__B net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11351_ _04482_ _07678_ vssd1 vssd1 vccd1 vccd1 _07680_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10274__C net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10302_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[18\] net772 net759 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06642_ sky130_fd_sc_hd__a22o_1
X_14070_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[12\] _04226_ _04256_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[44\]
+ _04357_ vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11282_ _07088_ _07154_ _07579_ _07589_ vssd1 vssd1 vccd1 vccd1 _07622_ sky130_fd_sc_hd__or4bb_1
XANTENNA__13866__B net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13021_ net3038 net3019 net865 vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__mux2_1
XANTENNA__08728__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10233_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[9\] _04646_ net799 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06573_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12262__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11732__A1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08679__C net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10164_ net1157 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[10\] net971
+ vssd1 vssd1 vccd1 vccd1 _06504_ sky130_fd_sc_hd__and3_1
XANTENNA__09137__A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input44_A wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1002 net1003 vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1013 net1014 vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__clkbuf_2
Xfanout1024 net1030 vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__buf_2
Xfanout1035 team_01_WB.instance_to_wrap.cpu.RU0.InstrRead vssd1 vssd1 vccd1 vccd1
+ net1035 sky130_fd_sc_hd__buf_2
Xfanout1046 net1049 vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__clkbuf_4
X_10095_ _06431_ _06432_ _06433_ _06434_ vssd1 vssd1 vccd1 vccd1 _06435_ sky130_fd_sc_hd__or4_1
Xfanout1057 net1058 vssd1 vssd1 vccd1 vccd1 net1057 sky130_fd_sc_hd__clkbuf_2
X_17760_ clknet_leaf_117_wb_clk_i _03436_ _01700_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14972_ net1249 vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__inv_2
XANTENNA__08976__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1068 team_01_WB.instance_to_wrap.cpu.f0.i\[27\] vssd1 vssd1 vccd1 vccd1 net1068
+ sky130_fd_sc_hd__clkbuf_4
Xfanout1079 net1080 vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__clkbuf_2
X_13923_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[14\] _04215_ net572 vssd1
+ vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__a21boi_1
X_16711_ clknet_leaf_107_wb_clk_i _02398_ _00694_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17691_ clknet_leaf_128_wb_clk_i _03375_ _01632_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11606__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08361__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16642_ clknet_leaf_55_wb_clk_i _02329_ _00625_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13854_ net1180 net1067 net1701 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[15\]
+ sky130_fd_sc_hd__and3b_1
X_12805_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] net1062 net364 _03631_
+ vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__a22o_1
X_16573_ clknet_leaf_68_wb_clk_i _02260_ _00556_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_13785_ _04156_ _01836_ vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__nand2_1
XANTENNA__09303__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10997_ net368 _07325_ _07336_ net552 _07335_ vssd1 vssd1 vccd1 vccd1 _07337_ sky130_fd_sc_hd__o221a_1
XFILLER_0_123_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15524_ net1222 vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__inv_2
XANTENNA__10449__C net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12736_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] net1061 net362 _03584_
+ vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_26_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09861__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10471__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15455_ net1312 vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__inv_2
X_12667_ net2215 net237 net387 vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__mux2_1
XANTENNA__12437__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12748__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14406_ net1361 vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11618_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[28\] _07088_ net715 vssd1 vssd1
+ vccd1 vccd1 _07832_ sky130_fd_sc_hd__mux2_1
XANTENNA__09613__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15386_ net1373 vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__inv_2
X_12598_ net2489 net200 net395 vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17125_ clknet_leaf_50_wb_clk_i _02812_ _01108_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11420__A0 team_01_WB.instance_to_wrap.cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_25_466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08967__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17913__1444 vssd1 vssd1 vccd1 vccd1 _17913__1444/HI net1444 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_133_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14337_ net1330 vssd1 vssd1 vccd1 vccd1 _00131_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11549_ net1577 net1173 vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold507 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2042 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold518 team_01_WB.instance_to_wrap.a1.ADR_I\[16\] vssd1 vssd1 vccd1 vccd1 net2053
+ sky130_fd_sc_hd__dlygate4sd3_1
X_17056_ clknet_leaf_48_wb_clk_i _02743_ _01039_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold529 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2064 sky130_fd_sc_hd__dlygate4sd3_1
X_14268_ net1225 vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16007_ net1357 vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__inv_2
X_13219_ net3092 net353 net349 team_01_WB.instance_to_wrap.cpu.f0.i\[31\] vssd1 vssd1
+ vccd1 vccd1 _01931_ sky130_fd_sc_hd__a22o_1
XANTENNA__12172__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13712__A2 _04504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14199_ _04156_ _01836_ _04181_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12025__X _07954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10526__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12920__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14888__A net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1207 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2742 sky130_fd_sc_hd__dlygate4sd3_1
X_08760_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[4\] net646 _05077_ _05080_
+ _05091_ vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_29_Left_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1218 team_01_WB.instance_to_wrap.cpu.f0.state\[0\] vssd1 vssd1 vccd1 vccd1 net2753
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17958_ net1473 vssd1 vssd1 vccd1 vccd1 la_data_out[0] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_81_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold1229 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2764 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09144__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16909_ clknet_leaf_67_wb_clk_i _02596_ _00892_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_08691_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[7\] net670 _05012_ _05018_
+ _05020_ vssd1 vssd1 vccd1 vccd1 _05031_ sky130_fd_sc_hd__a2111o_1
X_17889_ net107 vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_10_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_109_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11516__S team_01_WB.instance_to_wrap.cpu.DM0.next_enable vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08352__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13228__B2 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09213__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09312_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[22\] net684 _05632_
+ _05634_ _05635_ vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_24_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09243_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[21\] net678 net662 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__a22o_1
XANTENNA__12347__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_38_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout231_A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12739__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09174_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[16\] net656 _05511_
+ _05512_ _05513_ vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13400__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08958__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08125_ _04472_ team_01_WB.instance_to_wrap.cpu.f0.num\[23\] team_01_WB.instance_to_wrap.cpu.f0.num\[19\]
+ _04475_ vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16116__Q team_01_WB.instance_to_wrap.cpu.f0.data_adr\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1140_A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10765__A2 _05898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08056_ _04530_ _04531_ _04533_ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__or3_1
XFILLER_0_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09883__C net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13164__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12082__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1026_X net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1405_A net1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10517__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09383__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11190__A2 _07526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout486_X net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08958_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[6\] net666 _05268_ _05270_
+ _05287_ vssd1 vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_129_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08889_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[2\] net936 vssd1
+ vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout653_X net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10920_ net370 _07257_ _07259_ net336 _07258_ vssd1 vssd1 vccd1 vccd1 _07260_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout820_X net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10851_ _06601_ _07189_ _06532_ _06594_ vssd1 vssd1 vccd1 vccd1 _07191_ sky130_fd_sc_hd__a211oi_2
XANTENNA__09123__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout918_X net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10269__C net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13570_ net720 _07251_ net1073 vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09843__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10782_ net554 _07121_ vssd1 vssd1 vccd1 vccd1 _07122_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12521_ net2290 net288 net408 vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12257__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15240_ net1376 vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__inv_2
X_12452_ net3009 net308 net418 vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__mux2_1
X_11403_ _04471_ _07713_ vssd1 vssd1 vccd1 vccd1 _07725_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_10_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15171_ net1249 vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12383_ net2869 net299 net425 vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14122_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[14\] _04226_ _04252_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[110\]
+ _04407_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_91_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11334_ _07665_ net1817 _07655_ vssd1 vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13155__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13088__S net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14053_ _04224_ _04238_ vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__nor2_1
X_11265_ _06922_ _06930_ _07071_ _07603_ _07604_ vssd1 vssd1 vccd1 vccd1 _07605_ sky130_fd_sc_hd__a32o_1
XFILLER_0_120_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10508__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13004_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[82\] net2952 net863 vssd1 vssd1
+ vccd1 vccd1 _02121_ sky130_fd_sc_hd__mux2_1
X_10216_ _06534_ _06553_ _06554_ _06555_ vssd1 vssd1 vccd1 vccd1 _06556_ sky130_fd_sc_hd__or4_1
XANTENNA__09374__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11196_ net333 net336 _07362_ vssd1 vssd1 vccd1 vccd1 _07536_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17812_ clknet_leaf_91_wb_clk_i _03488_ _01752_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[82\]
+ sky130_fd_sc_hd__dfrtp_1
X_10147_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[11\] net817 net738 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[11\]
+ _06474_ vssd1 vssd1 vccd1 vccd1 _06487_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_89_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14955_ net1396 vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__inv_2
X_17743_ clknet_leaf_98_wb_clk_i _03419_ _01683_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[13\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_89_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10078_ net1138 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[7\] net958 vssd1
+ vssd1 vccd1 vccd1 _06418_ sky130_fd_sc_hd__and3_1
X_13906_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[7\] _04204_ _04205_ vssd1
+ vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__o21a_1
X_17674_ clknet_leaf_157_wb_clk_i _03359_ _01615_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10141__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14886_ net1400 vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__inv_2
XANTENNA__10692__A1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13837_ net2427 net830 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[30\]
+ sky130_fd_sc_hd__and2_1
X_16625_ clknet_leaf_113_wb_clk_i _02312_ _00608_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13615__D1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15332__A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16556_ clknet_leaf_159_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[22\]
+ _00539_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13768_ net1184 _04155_ vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09834__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12719_ net2094 net289 net384 vssd1 vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__mux2_1
X_15507_ net1419 vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16487_ clknet_leaf_156_wb_clk_i _02241_ _00470_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12167__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13699_ net1816 _04106_ _04120_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[10\]
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_100_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10995__A2 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15438_ net1294 vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_80_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11859__X _07948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15369_ net1295 vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__inv_2
Xhold304 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1839 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17108_ clknet_leaf_22_wb_clk_i _02795_ _01091_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold315 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1850 sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[29\] vssd1 vssd1 vccd1 vccd1 net1861
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[1\] vssd1 vssd1 vccd1 vccd1
+ net1872 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13146__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold348 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1883 sky130_fd_sc_hd__dlygate4sd3_1
X_09930_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[4\] net741 net771 vssd1
+ vssd1 vccd1 vccd1 _06270_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17039_ clknet_leaf_37_wb_clk_i _02726_ _01022_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold359 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1894 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout806 _04641_ vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__buf_6
X_09861_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[12\] net820 net783 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06201_ sky130_fd_sc_hd__a22o_1
Xfanout817 net818 vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__buf_6
Xfanout828 _04578_ vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__buf_2
XANTENNA__09208__C net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout839 _03734_ vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__buf_2
XANTENNA__11172__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08812_ net602 _05150_ _05116_ vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__a21o_1
XANTENNA__12630__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13449__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09792_ net374 _06131_ vssd1 vssd1 vccd1 vccd1 _06132_ sky130_fd_sc_hd__nand2_1
Xhold1004 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2539 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1015 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2550 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10380__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1026 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2561 sky130_fd_sc_hd__dlygate4sd3_1
X_08743_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[4\] net919 vssd1
+ vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__and3_1
Xhold1037 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[16\] vssd1 vssd1 vccd1 vccd1
+ net2572 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09505__A net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1048 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[58\] vssd1 vssd1 vccd1 vccd1
+ net2594 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout279_A _07917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08674_ net1006 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[7\] net900 vssd1
+ vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_124_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13606__D1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1090_A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout446_A _07959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1188_A net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_46_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08408__X _04748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13621__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08782__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12077__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout613_A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout234_X net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1355_A net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09226_ net597 _05564_ _05565_ vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_1_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13968__Y _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09157_ net1017 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[16\] net893
+ vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout401_X net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1143_X net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08108_ _04504_ net1176 vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__and2_1
X_09088_ net1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[13\] net930
+ vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout982_A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13137__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08039_ net1674 net567 net345 team_01_WB.instance_to_wrap.cpu.f0.i\[16\] vssd1 vssd1
+ vccd1 vccd1 _03552_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_55_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold860 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2395 sky130_fd_sc_hd__dlygate4sd3_1
Xhold871 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2406 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08303__B net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1408_X net1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold882 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2417 sky130_fd_sc_hd__dlygate4sd3_1
Xhold893 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2428 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11050_ net517 _06339_ vssd1 vssd1 vccd1 vccd1 _07390_ sky130_fd_sc_hd__nand2_1
XANTENNA__09356__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout770_X net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09118__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout868_X net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10001_ net552 net541 net561 vssd1 vssd1 vccd1 vccd1 _06341_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12540__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10371__B1 _05566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09108__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14101__A2 _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14040__B net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1560 team_01_WB.instance_to_wrap.cpu.K0.code\[2\] vssd1 vssd1 vccd1 vccd1 net3095
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1571 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net3106 sky130_fd_sc_hd__dlygate4sd3_1
X_14740_ net1197 vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__inv_2
X_11952_ net2054 net295 net477 vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17912__1443 vssd1 vssd1 vccd1 vccd1 _17912__1443/HI net1443 sky130_fd_sc_hd__conb_1
Xhold1582 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[18\] vssd1 vssd1 vccd1 vccd1
+ net3117 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_28_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1593 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net3128 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10903_ _04883_ _06672_ vssd1 vssd1 vccd1 vccd1 _07243_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14671_ net1225 vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_64_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11883_ net1986 net300 net483 vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_84_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12776__A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16410_ clknet_leaf_123_wb_clk_i _02164_ _00393_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13622_ net720 _07531_ net1076 vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__o21a_1
X_10834_ _06194_ _07173_ _06599_ _06164_ vssd1 vssd1 vccd1 vccd1 _07174_ sky130_fd_sc_hd__o211a_1
X_17390_ clknet_leaf_27_wb_clk_i _03077_ _01373_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16525__CLK clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11623__A0 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16341_ clknet_leaf_122_wb_clk_i _02095_ _00324_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[64\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13553_ net185 _04002_ _04003_ net723 vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__a211o_1
X_17909__1520 vssd1 vssd1 vccd1 vccd1 net1520 _17909__1520/LO sky130_fd_sc_hd__conb_1
X_10765_ _04706_ net513 _05898_ net504 net548 net537 vssd1 vssd1 vccd1 vccd1 _07105_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_137_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10977__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12504_ net3105 net265 net407 vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__mux2_1
X_16272_ clknet_leaf_88_wb_clk_i _00000_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13484_ _03848_ _03944_ vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10696_ _06936_ _06943_ net535 vssd1 vssd1 vccd1 vccd1 _07036_ sky130_fd_sc_hd__mux2_1
X_18011_ net1510 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__buf_2
X_15223_ net1244 vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12435_ net2049 net271 net417 vssd1 vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__mux2_1
XANTENNA__12715__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15154_ net1290 vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09595__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_73_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12366_ net1863 net203 net423 vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_136_Right_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13128__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14105_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[37\] _04221_ _04260_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[61\]
+ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11317_ team_01_WB.instance_to_wrap.cpu.f0.state\[5\] _04506_ team_01_WB.instance_to_wrap.cpu.f0.state\[8\]
+ _04524_ _00019_ vssd1 vssd1 vccd1 vccd1 _07654_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_39_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15085_ net1264 vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__inv_2
X_12297_ net1935 net246 net433 vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__mux2_1
X_14036_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[58\] _04260_ _04266_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[18\]
+ _04313_ vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__a221o_1
XANTENNA_output75_A net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09347__A2 _04776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11248_ _07555_ _07580_ _07586_ _07587_ vssd1 vssd1 vccd1 vccd1 _07588_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_56_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08555__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12450__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10362__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11179_ net338 _07065_ _07518_ vssd1 vssd1 vccd1 vccd1 _07519_ sky130_fd_sc_hd__a21o_1
XANTENNA__08867__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15987_ net1368 vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17726_ clknet_leaf_150_wb_clk_i _03403_ _01667_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__10114__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14938_ net1370 vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__inv_2
X_17657_ clknet_leaf_2_wb_clk_i _03342_ _01598_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14869_ net1282 vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_102_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15062__A net1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11590__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16608_ clknet_leaf_45_wb_clk_i _02295_ _00591_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_08390_ _04708_ _04717_ _04726_ net710 vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__nor4_1
XANTENNA__09807__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17588_ clknet_leaf_130_wb_clk_i _03275_ _01547_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.code\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13603__A1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09698__C net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_154_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16539_ clknet_leaf_6_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[5\]
+ _00522_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11090__A1 _04706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09011_ net1021 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[9\] net936 vssd1
+ vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12625__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13310__A team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_79_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold101 net124 vssd1 vssd1 vccd1 vccd1 net1636 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09586__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold112 net114 vssd1 vssd1 vccd1 vccd1 net1647 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 net81 vssd1 vssd1 vccd1 vccd1 net1658 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08404__A _04743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold134 team_01_WB.instance_to_wrap.cpu.f0.write_data\[8\] vssd1 vssd1 vccd1 vccd1
+ net1669 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold145 team_01_WB.instance_to_wrap.cpu.f0.write_data\[15\] vssd1 vssd1 vccd1 vccd1
+ net1680 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 team_01_WB.instance_to_wrap.a1.ADR_I\[22\] vssd1 vssd1 vccd1 vccd1 net1691
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 net132 vssd1 vssd1 vccd1 vccd1 net1702 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold178 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[7\] vssd1 vssd1 vccd1 vccd1
+ net1713 sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ _05076_ _06252_ vssd1 vssd1 vccd1 vccd1 _06253_ sky130_fd_sc_hd__xor2_1
XANTENNA__09338__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold189 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 net1724
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout603 _04754_ vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__buf_4
Xfanout614 _07636_ vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout396_A _03567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout625 net627 vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__buf_4
Xfanout636 net637 vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__clkbuf_2
X_09844_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[13\] net787 net760 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06184_ sky130_fd_sc_hd__a22o_1
XANTENNA__12360__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout647 _04825_ vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__buf_2
Xfanout658 _04813_ vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__buf_6
XANTENNA_fanout1103_A net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout669 net670 vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__buf_6
XANTENNA__08777__C net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09775_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[15\] net789 net775 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_126_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08726_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[5\] net660 _05044_ _05047_
+ _05052_ vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10105__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08849__A1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08657_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[10\] net666 _04972_
+ _04974_ _04985_ vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10656__B2 _06906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout730_A net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1093_X net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout449_X net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11704__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08588_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[15\] net668 net655 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12883__X _03663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout616_X net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10550_ _06888_ _06889_ net538 vssd1 vssd1 vccd1 vccd1 _06890_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09209_ net1083 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[17\] net926
+ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__and3_1
X_10481_ _06781_ _06815_ vssd1 vssd1 vccd1 vccd1 _06821_ sky130_fd_sc_hd__nor2_1
XANTENNA__12535__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12220_ net2141 net317 net446 vssd1 vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_920 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09577__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08314__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10563__B _06902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout985_X net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12151_ net1719 net294 net453 vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__mux2_1
XANTENNA__10592__B1 _06906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11102_ net555 net332 _07396_ net337 net370 vssd1 vssd1 vccd1 vccd1 _07442_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_4_5__f_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09329__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12082_ net2227 net300 net459 vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__mux2_1
Xhold690 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2225 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13530__B1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15910_ net1415 vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__inv_2
X_11033_ _07368_ _07371_ _07372_ vssd1 vssd1 vccd1 vccd1 _07373_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_34_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12270__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16890_ clknet_leaf_82_wb_clk_i _02577_ _00873_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08687__C net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15841_ net1326 vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_138_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_138_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_51_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15772_ net1217 vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__inv_2
X_12984_ net2858 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[110\] net855 vssd1 vssd1
+ vccd1 vccd1 _02141_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1390 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2925 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_82_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17511_ clknet_leaf_100_wb_clk_i _03198_ _01494_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_26_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14723_ net1196 vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__inv_2
X_11935_ net2298 net201 net475 vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__mux2_1
X_17442_ clknet_leaf_56_wb_clk_i _03129_ _01425_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_14654_ net1238 vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__inv_2
X_11866_ net2699 net206 net485 vssd1 vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13605_ _04029_ _04046_ vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__nor2_1
X_10817_ net512 _05963_ _06779_ _06811_ net548 net533 vssd1 vssd1 vccd1 vccd1 _07157_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_131_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17373_ clknet_leaf_64_wb_clk_i _03060_ _01356_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_14585_ net1413 vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__inv_2
X_11797_ net3032 net247 net493 vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13536_ net986 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] _03988_ _03989_
+ vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__a22o_1
X_16324_ clknet_leaf_120_wb_clk_i net2603 _00307_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[47\]
+ sky130_fd_sc_hd__dfrtp_1
X_10748_ net563 _06825_ _07057_ _07087_ vssd1 vssd1 vccd1 vccd1 _07088_ sky130_fd_sc_hd__a31o_2
XFILLER_0_55_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16255_ clknet_leaf_152_wb_clk_i net1546 _00243_ vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12445__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13467_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] _05655_ vssd1 vssd1
+ vccd1 vccd1 _03928_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10679_ net563 _06829_ _06962_ _07018_ vssd1 vssd1 vccd1 vccd1 _07019_ sky130_fd_sc_hd__a31o_2
XANTENNA__10754__A _04844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14226__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15206_ net1404 vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__inv_2
X_12418_ net2472 net311 net419 vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__mux2_1
X_16186_ clknet_leaf_1_wb_clk_i _01946_ _00174_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13398_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] _05495_ vssd1 vssd1
+ vccd1 vccd1 _03859_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_58_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15137_ net1279 vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__inv_2
X_12349_ net1892 net279 net428 vssd1 vssd1 vccd1 vccd1 _02646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15068_ net1246 vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_147_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14019_ net1561 net605 _04309_ net1183 vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__o211a_1
XANTENNA__11585__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12180__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_65_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10886__A1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09560_ _05760_ _05781_ vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__xnor2_1
X_08511_ net1081 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[18\] net914
+ vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_19_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17709_ clknet_leaf_134_wb_clk_i _03393_ _01650_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[30\]
+ sky130_fd_sc_hd__dfrtp_4
X_09491_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[30\] net695 net674 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[30\]
+ _05821_ vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_121_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08442_ net1117 net1120 net1123 net1126 vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__and4_1
XFILLER_0_93_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08373_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__or2_2
XFILLER_0_18_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout311_A _07931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12355__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1053_A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout409_A _03564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17911__1442 vssd1 vssd1 vccd1 vccd1 _17911__1442/HI net1442 sky130_fd_sc_hd__conb_1
XANTENNA__16124__Q team_01_WB.instance_to_wrap.cpu.f0.data_adr\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1220_A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1318_A net1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09891__C net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout680_A _04787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout400 _03566_ vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__buf_4
Xfanout1409 net1428 vssd1 vssd1 vccd1 vccd1 net1409 sky130_fd_sc_hd__buf_2
Xfanout411 _03563_ vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__buf_6
XANTENNA_fanout778_A _04666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout399_X net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout422 _03561_ vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__buf_6
XANTENNA__12090__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout433 _07964_ vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__buf_6
Xfanout444 _07959_ vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout455 _07956_ vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__buf_6
XANTENNA_fanout1106_X net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout466 _07954_ vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09827_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[13\] net779 net777 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[13\]
+ _06166_ vssd1 vssd1 vccd1 vccd1 _06167_ sky130_fd_sc_hd__a221o_1
Xfanout477 _07950_ vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__buf_6
Xfanout488 _07947_ vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout566_X net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout499 net502 vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__buf_6
XANTENNA_fanout945_A net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09758_ net582 _06097_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] net627
+ vssd1 vssd1 vccd1 vccd1 _06098_ sky130_fd_sc_hd__a2bb2o_2
X_08709_ net1098 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[5\] net913 vssd1
+ vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout733_X net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09689_ _06025_ _06026_ _06027_ _06028_ vssd1 vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__or4_1
XANTENNA__10398__X _06738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11720_ net714 _07308_ vssd1 vssd1 vccd1 vccd1 _07913_ sky130_fd_sc_hd__nand2_1
XANTENNA__10558__B _05151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout900_X net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11651_ net2218 net201 net499 vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__mux2_1
XANTENNA__09131__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10277__C net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10602_ net550 _06526_ vssd1 vssd1 vccd1 vccd1 _06942_ sky130_fd_sc_hd__nor2_1
XANTENNA__09798__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14370_ net1208 vssd1 vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11582_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] _07798_ vssd1 vssd1 vccd1
+ vccd1 _07799_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08970__C net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13321_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[20\] net826 _03799_ _03800_
+ vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10533_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[31\] net656 net705 vssd1
+ vssd1 vccd1 vccd1 _06873_ sky130_fd_sc_hd__a21o_1
XANTENNA__12265__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16040_ clknet_leaf_88_wb_clk_i _01834_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13252_ net610 _07710_ net1069 vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__a21o_1
XANTENNA_input74_A wbs_we_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11389__B _07696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10464_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[26\] net757 _06789_ _06790_
+ _06792_ vssd1 vssd1 vccd1 vccd1 _06804_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_20_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12203_ net2118 net240 net443 vssd1 vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__mux2_1
X_13183_ net1177 net837 team_01_WB.instance_to_wrap.a1.prev_BUSY_O vssd1 vssd1 vccd1
+ vccd1 _03739_ sky130_fd_sc_hd__or3b_1
X_10395_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[16\] net819 net777 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06735_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12134_ net3002 net200 net451 vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09970__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17991_ net635 vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10580__Y _06920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16942_ clknet_leaf_38_wb_clk_i _02629_ _00925_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_12065_ net2264 net208 net461 vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11016_ _05618_ net507 vssd1 vssd1 vccd1 vccd1 _07356_ sky130_fd_sc_hd__xor2_1
XANTENNA__09722__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16873_ clknet_leaf_39_wb_clk_i _02560_ _00856_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15824_ net1202 vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_149_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_126_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09603__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15755_ net1342 vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__inv_2
X_12967_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[119\] net1888 net856 vssd1 vssd1
+ vccd1 vccd1 _02158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11918_ net2954 net298 net481 vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__mux2_1
X_14706_ net1193 vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15686_ net1384 vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__inv_2
X_12898_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[23\] net1036 vssd1 vssd1 vccd1
+ vccd1 _03674_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17425_ clknet_leaf_113_wb_clk_i _03112_ _01408_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11849_ net2644 net281 net488 vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__mux2_1
XANTENNA__12883__B1_N net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14637_ net1270 vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17356_ clknet_leaf_147_wb_clk_i _03043_ _01339_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_14568_ net1352 vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_35_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_28_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12793__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16307_ clknet_leaf_116_wb_clk_i _02061_ _00290_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12175__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13519_ net988 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] _03974_ _03975_
+ vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__a22o_1
XANTENNA__13990__B1 _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14499_ net1415 vssd1 vssd1 vccd1 vccd1 _00293_ sky130_fd_sc_hd__inv_2
X_17287_ clknet_leaf_107_wb_clk_i _02974_ _01270_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload10 clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload10/Y sky130_fd_sc_hd__clkinv_4
Xclkload21 clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload21/Y sky130_fd_sc_hd__bufinv_16
X_16238_ clknet_leaf_152_wb_clk_i net1621 _00226_ vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__dfrtp_1
Xclkload32 clknet_leaf_153_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload32/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_70_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload43 clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload43/X sky130_fd_sc_hd__clkbuf_8
Xclkload54 clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload54/Y sky130_fd_sc_hd__bufinv_16
Xclkload65 clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload65/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_149_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload76 clknet_leaf_59_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload76/Y sky130_fd_sc_hd__inv_6
XANTENNA__10771__X _07111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16169_ clknet_leaf_3_wb_clk_i _00011_ _00157_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
Xclkload87 clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload87/Y sky130_fd_sc_hd__inv_6
XANTENNA__08889__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload98 clknet_leaf_130_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload98/Y sky130_fd_sc_hd__inv_6
XFILLER_0_62_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10020__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08991_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[8\] net671 _05328_ _05329_
+ _05330_ vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__09961__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Left_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10859__A1 _06707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09713__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_4__f_wb_clk_i_X clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09612_ _05949_ _05950_ _05951_ vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__or3_1
XFILLER_0_92_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09543_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[28\] net746 _05872_ _05874_
+ _05881_ vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11462__B1_N net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout261_A _07880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout359_A _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10087__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09474_ net1083 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[30\] net891
+ vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17929__1446 vssd1 vssd1 vccd1 vccd1 _17929__1446/HI net1446 sky130_fd_sc_hd__conb_1
XANTENNA__16119__Q team_01_WB.instance_to_wrap.cpu.f0.data_adr\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08425_ net1119 net1122 net1125 net1116 vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_149_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout526_A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1268_A net1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08356_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[30\] net782 net755 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09886__C net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08790__C net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload4 clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload4/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__12784__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12085__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08287_ _04625_ _04626_ vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__nor2_1
XANTENNA__10795__B1 _07134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11002__B net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10547__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1223_X net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10011__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10180_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[10\] net788 net754 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06520_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout683_X net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1206 net1207 vssd1 vssd1 vccd1 vccd1 net1206 sky130_fd_sc_hd__buf_4
Xfanout1217 net1219 vssd1 vssd1 vccd1 vccd1 net1217 sky130_fd_sc_hd__buf_4
Xfanout1228 net1229 vssd1 vssd1 vccd1 vccd1 net1228 sky130_fd_sc_hd__buf_2
Xfanout230 net232 vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08311__B net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout241 net244 vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__buf_2
XANTENNA__09165__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1239 net1241 vssd1 vssd1 vccd1 vccd1 net1239 sky130_fd_sc_hd__buf_2
Xfanout252 _07904_ vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11282__C_N _07579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout263 _07880_ vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__buf_2
XANTENNA_fanout850_X net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17993__1505 vssd1 vssd1 vccd1 vccd1 _17993__1505/HI net1505 sky130_fd_sc_hd__conb_1
XANTENNA__09126__C net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout274 net275 vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__clkbuf_2
Xfanout285 _07896_ vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__buf_1
XANTENNA_fanout948_X net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout296 net297 vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__clkbuf_2
X_13870_ net1177 net1064 net1615 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[31\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_119_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08965__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12821_ net1569 net640 net608 _03643_ vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__a22o_1
XANTENNA__09468__A1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12752_ net364 _03594_ _03595_ net1062 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__a32o_1
XFILLER_0_57_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15540_ net1380 vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11703_ net612 _07806_ _07899_ _07898_ vssd1 vssd1 vccd1 vccd1 _07900_ sky130_fd_sc_hd__a31o_1
X_15471_ net1299 vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__inv_2
X_12683_ net2068 net305 net390 vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__mux2_1
XANTENNA__08691__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17210_ clknet_leaf_79_wb_clk_i _02897_ _01193_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_14422_ net1310 vssd1 vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__inv_2
X_11634_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] _07817_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\]
+ vssd1 vssd1 vccd1 vccd1 _07845_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_46_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08326__X _04666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14353_ net1333 vssd1 vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__inv_2
X_17141_ clknet_leaf_111_wb_clk_i _02828_ _01124_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11565_ net3142 net155 team_01_WB.instance_to_wrap.cpu.K0.next_state vssd1 vssd1
+ vccd1 vccd1 _03274_ sky130_fd_sc_hd__mux2_1
XANTENNA__10786__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13304_ _07686_ _07711_ _03786_ net587 vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_42_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10516_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[31\] net764 net622 vssd1
+ vssd1 vccd1 vccd1 _06856_ sky130_fd_sc_hd__o21a_1
X_17072_ clknet_leaf_147_wb_clk_i _02759_ _01055_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14284_ net1336 vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__inv_2
X_11496_ net367 _07775_ net2001 net875 vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_150_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13235_ net3035 net355 net351 team_01_WB.instance_to_wrap.cpu.f0.i\[15\] vssd1 vssd1
+ vccd1 vccd1 _01915_ sky130_fd_sc_hd__a22o_1
X_16023_ net1327 vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_94_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10447_ net1147 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[26\] _04660_
+ vssd1 vssd1 vccd1 vccd1 _06787_ sky130_fd_sc_hd__and3_1
XANTENNA__10538__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13166_ net1915 net847 net839 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[10\] vssd1
+ vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__a22o_1
X_10378_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[16\] net811 net739 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[16\]
+ _06716_ vssd1 vssd1 vccd1 vccd1 _06718_ sky130_fd_sc_hd__a221o_1
X_12117_ net2291 net296 net458 vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_153_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_153_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_17974_ net1489 vssd1 vssd1 vccd1 vccd1 la_data_out[16] sky130_fd_sc_hd__buf_2
X_13097_ net70 net69 net41 net40 vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__or4_1
XFILLER_0_97_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12048_ net2113 net282 net466 vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__mux2_1
X_16925_ clknet_leaf_69_wb_clk_i _02612_ _00908_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11502__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15335__A net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16856_ clknet_leaf_50_wb_clk_i _02543_ _00839_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_15807_ net1200 vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__inv_2
X_16787_ clknet_leaf_22_wb_clk_i _02474_ _00770_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13999_ _04238_ _04242_ vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11266__A1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15738_ net1372 vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15669_ net1277 vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08210_ net2712 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[63\] net1048 vssd1 vssd1
+ vccd1 vccd1 _03477_ sky130_fd_sc_hd__mux2_1
XANTENNA__11802__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17408_ clknet_leaf_48_wb_clk_i _03095_ _01391_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_09190_ net1163 net620 net593 vssd1 vssd1 vccd1 vccd1 _05530_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10926__B _07227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08141_ _04472_ team_01_WB.instance_to_wrap.cpu.f0.num\[23\] team_01_WB.instance_to_wrap.cpu.f0.num\[20\]
+ _04474_ _04593_ vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__a221o_1
X_17339_ clknet_leaf_71_wb_clk_i _03026_ _01322_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10777__A0 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10241__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08072_ team_01_WB.instance_to_wrap.cpu.f0.i\[5\] _04524_ vssd1 vssd1 vccd1 vccd1
+ _04549_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload110 clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload110/Y sky130_fd_sc_hd__clkinv_8
Xclkload121 clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload121/Y sky130_fd_sc_hd__clkinv_4
Xclkload132 clknet_leaf_82_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload132/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_31_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload143 clknet_leaf_84_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload143/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_113_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12633__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10529__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09395__B1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09934__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11757__B team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08412__A _04708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10544__A3 _05835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08974_ net1087 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[8\] net914 vssd1
+ vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__and3_1
XANTENNA__09227__B _05566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1016_A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold16 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[1\] vssd1 vssd1 vccd1 vccd1
+ net1551 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold27 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[5\] vssd1 vssd1 vccd1 vccd1 net1562
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14140__B1 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold38 net95 vssd1 vssd1 vccd1 vccd1 net1573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 team_01_WB.instance_to_wrap.cpu.f0.write_data\[27\] vssd1 vssd1 vccd1 vccd1
+ net1584 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout476_A _07950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08785__C net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1385_A net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09526_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[29\] net765 net624 vssd1
+ vssd1 vccd1 vccd1 _05866_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_149_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09457_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[29\] net692 net660 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout431_X net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout908_A net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout529_X net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08408_ _04738_ _04746_ vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09388_ net601 _05727_ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08339_ net1131 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[30\] net965
+ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__and3_1
XFILLER_0_85_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08306__B net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10232__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11350_ _04482_ _07678_ vssd1 vssd1 vccd1 vccd1 _07679_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout898_X net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10301_ _06639_ _06640_ vssd1 vssd1 vccd1 vccd1 _06641_ sky130_fd_sc_hd__nand2_1
X_11281_ net562 _07612_ _07613_ _07620_ vssd1 vssd1 vccd1 vccd1 _07621_ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12543__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13020_ net2779 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[74\] net863 vssd1 vssd1
+ vccd1 vccd1 _02105_ sky130_fd_sc_hd__mux2_1
XANTENNA__09386__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10232_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[9\] net808 net736 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[9\]
+ _06570_ vssd1 vssd1 vccd1 vccd1 _06572_ sky130_fd_sc_hd__a221o_1
XANTENNA__09925__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_1_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11732__A2 _07507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10163_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[10\] net792 net778 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06503_ sky130_fd_sc_hd__a22o_1
Xfanout1003 net1015 vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__clkbuf_4
Xfanout1014 net1015 vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10290__C net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1025 net1026 vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__clkbuf_2
Xfanout1036 net1037 vssd1 vssd1 vccd1 vccd1 net1036 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input37_A gpio_in[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1047 net1048 vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__clkbuf_4
X_10094_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[7\] net801 net749 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06434_ sky130_fd_sc_hd__a22o_1
X_14971_ net1254 vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__inv_2
Xfanout1058 net1059 vssd1 vssd1 vccd1 vccd1 net1058 sky130_fd_sc_hd__buf_2
Xfanout1069 team_01_WB.instance_to_wrap.cpu.f0.i\[22\] vssd1 vssd1 vccd1 vccd1 net1069
+ sky130_fd_sc_hd__clkbuf_4
X_16710_ clknet_leaf_73_wb_clk_i _02397_ _00693_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13922_ _04215_ net571 _04214_ vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__and3b_1
XFILLER_0_156_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17690_ clknet_leaf_127_wb_clk_i _03374_ _01631_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_107_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16641_ clknet_leaf_55_wb_clk_i _02328_ _00624_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13853_ net1180 net1067 net3175 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[14\]
+ sky130_fd_sc_hd__and3b_1
XANTENNA__10299__A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12804_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[8\] _07290_ net1035 vssd1 vssd1
+ vccd1 vccd1 _03631_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16572_ clknet_leaf_64_wb_clk_i _02259_ _00555_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_13784_ _04162_ _04164_ vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__xnor2_1
X_10996_ _06398_ net334 net332 vssd1 vssd1 vccd1 vccd1 _07336_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09440__X _05780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15523_ net1222 vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__inv_2
X_12735_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[30\] _07019_ net1032 vssd1 vssd1
+ vccd1 vccd1 _03584_ sky130_fd_sc_hd__mux2_1
XANTENNA__12718__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11622__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10471__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12666_ net2981 net269 net387 vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__mux2_1
X_15454_ net1350 vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12748__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14405_ net1361 vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__inv_2
X_11617_ net2703 net218 net501 vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15385_ net1231 vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12597_ net2093 net203 net395 vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17124_ clknet_leaf_73_wb_clk_i _02811_ _01107_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_14336_ net1338 vssd1 vssd1 vccd1 vccd1 _00130_ sky130_fd_sc_hd__inv_2
X_11548_ net1552 net1173 vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__and2_1
XFILLER_0_135_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold508 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2043 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12453__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17055_ clknet_leaf_41_wb_clk_i _02742_ _01038_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold519 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2054 sky130_fd_sc_hd__dlygate4sd3_1
X_14267_ net1224 vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__inv_2
X_11479_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[23\] net579 vssd1 vssd1 vccd1
+ vccd1 _07767_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11210__X _07550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13218_ team_01_WB.instance_to_wrap.cpu.f0.state\[6\] _03740_ vssd1 vssd1 vccd1 vccd1
+ _03742_ sky130_fd_sc_hd__nor2_1
X_16006_ net1331 vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__inv_2
XANTENNA__09377__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09916__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14198_ net1588 _04462_ _04463_ vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__o21a_1
XFILLER_0_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12920__A1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13149_ net1678 net850 net842 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[27\] vssd1
+ vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14122__B1 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17957_ net1472 vssd1 vssd1 vccd1 vccd1 irq[2] sky130_fd_sc_hd__buf_2
Xhold1208 team_01_WB.instance_to_wrap.cpu.f0.num\[29\] vssd1 vssd1 vccd1 vccd1 net2743
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1219 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2754 sky130_fd_sc_hd__dlygate4sd3_1
X_16908_ clknet_leaf_149_wb_clk_i _02595_ _00891_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_08690_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[7\] net661 _05008_ _05013_
+ _05026_ vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__a2111o_1
X_17888_ net107 vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_109_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16839_ clknet_leaf_106_wb_clk_i _02526_ _00822_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13633__C1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10002__A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_50_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_105_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09311_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[22\] net665 _05622_
+ _05625_ _05638_ vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_119_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12628__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08655__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09242_ net1098 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[21\] net909
+ net657 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[21\] vssd1 vssd1 vccd1
+ vccd1 _05582_ sky130_fd_sc_hd__a32o_1
XANTENNA__10462__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12739__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09173_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[16\] net922
+ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout224_A _07827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08124_ _04481_ team_01_WB.instance_to_wrap.cpu.f0.num\[13\] team_01_WB.instance_to_wrap.cpu.f0.num\[12\]
+ _04482_ vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__o22a_1
XANTENNA__10214__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12871__B net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10765__A3 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08055_ _04527_ _04532_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__nor2_1
XANTENNA__12363__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1133_A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09368__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1300_A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1019_X net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14113__B1 _04266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08957_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[6\] net698 _05271_ _05282_
+ net707 vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout760_A net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout381_X net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout479_X net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout858_A net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1506_A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[5\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08888_ net1025 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[2\] net902 vssd1
+ vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout646_X net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10850_ _06601_ _07189_ _06594_ vssd1 vssd1 vccd1 vccd1 _07190_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09701__A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09509_ net1150 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[29\] net955
+ vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout813_X net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12538__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10781_ net529 _06967_ _07120_ _07119_ vssd1 vssd1 vccd1 vccd1 _07121_ sky130_fd_sc_hd__a31o_1
XFILLER_0_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12520_ net2240 net314 net409 vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__mux2_1
XANTENNA__08317__A net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ net2913 net310 net415 vssd1 vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11402_ net323 _07723_ _07724_ vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__and3_1
XFILLER_0_151_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15170_ net1351 vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__inv_2
X_12382_ net2073 net277 net424 vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14121_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[94\] _04240_ _04268_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[78\]
+ vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11333_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[2\] team_01_WB.instance_to_wrap.cpu.f0.state\[4\]
+ _04555_ _07652_ vssd1 vssd1 vccd1 vccd1 _07665_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_91_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12273__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10582__A net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14054__A _04236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09359__B1 _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14052_ _04334_ _04336_ _04338_ _04340_ vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__or4_1
XFILLER_0_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11264_ net522 _07300_ net557 vssd1 vssd1 vccd1 vccd1 _07604_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13003_ net1542 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[91\] net861 vssd1 vssd1
+ vccd1 vccd1 _02122_ sky130_fd_sc_hd__mux2_1
X_10215_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[8\] net730 _06538_ _06542_
+ _06545_ vssd1 vssd1 vccd1 vccd1 _06555_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08031__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11195_ net327 _07534_ vssd1 vssd1 vccd1 vccd1 _07535_ sky130_fd_sc_hd__and2_1
X_17811_ clknet_leaf_94_wb_clk_i _03487_ _01751_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[81\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14104__B1 _04244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10146_ _06475_ _06478_ _06480_ _06485_ vssd1 vssd1 vccd1 vccd1 _06486_ sky130_fd_sc_hd__or4_1
XFILLER_0_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11617__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17742_ clknet_leaf_99_wb_clk_i _03418_ _01682_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[12\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_89_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10077_ net1138 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[7\] net973 vssd1
+ vssd1 vccd1 vccd1 _06417_ sky130_fd_sc_hd__and3_1
X_14954_ net1283 vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13905_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[7\] _04204_ net571 vssd1
+ vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__a21boi_1
X_17673_ clknet_leaf_0_wb_clk_i _03358_ _01614_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_14885_ net1287 vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload2_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16624_ clknet_leaf_144_wb_clk_i _02311_ _00607_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13836_ net1724 net830 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[29\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_76_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16555_ clknet_leaf_0_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[21\]
+ _00538_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12448__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13767_ team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[4\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[4\]
+ net604 vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__mux2_1
X_10979_ _06438_ net372 _06590_ _06562_ net550 net534 vssd1 vssd1 vccd1 vccd1 _07319_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_63_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15506_ net1291 vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12718_ net2580 net313 net385 vssd1 vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11641__B2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16486_ clknet_leaf_153_wb_clk_i _02240_ _00469_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_135_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13698_ team_01_WB.instance_to_wrap.cpu.c0.count\[10\] _04106_ _04119_ vssd1 vssd1
+ vccd1 vccd1 _04120_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_26_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16217__Q net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15437_ net1265 vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_80_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12649_ net2246 net309 net392 vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10195__C net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15368_ net1387 vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17107_ clknet_leaf_24_wb_clk_i _02794_ _01090_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12183__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14319_ net1358 vssd1 vssd1 vccd1 vccd1 _00113_ sky130_fd_sc_hd__inv_2
Xhold305 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold316 team_01_WB.instance_to_wrap.a1.ADR_I\[2\] vssd1 vssd1 vccd1 vccd1 net1851
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10492__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15299_ net1221 vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__inv_2
Xhold327 team_01_WB.instance_to_wrap.a1.ADR_I\[30\] vssd1 vssd1 vccd1 vccd1 net1862
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1873 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold349 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1884 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09058__A net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17038_ clknet_leaf_27_wb_clk_i _02725_ _01021_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout807 net810 vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__buf_6
X_09860_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[12\] net774 _06195_
+ _06199_ vssd1 vssd1 vccd1 vccd1 _06200_ sky130_fd_sc_hd__a211o_1
XANTENNA__12911__S net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout818 _04634_ vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__buf_6
Xfanout829 _04578_ vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__buf_2
X_08811_ net602 _05150_ _05116_ vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__a21oi_4
XANTENNA__09770__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09791_ _04947_ _06130_ vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1005 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2540 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2551 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1027 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2562 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08742_ net1012 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[4\] net897 vssd1
+ vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__and3_1
Xhold1038 _03422_ vssd1 vssd1 vccd1 vccd1 net2573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2584 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09522__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08673_ net1085 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[7\] net911 vssd1
+ vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__and3_1
XANTENNA__08876__A2 _04771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout341_A _06216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12358__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08628__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout439_A _07962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1083_A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire983_X net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10435__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09225_ net1163 net620 net593 net600 vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__a211o_1
XFILLER_0_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout606_A _03583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09156_ net1097 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[16\] net936
+ vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__and3_1
XANTENNA__07976__A team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11396__B1 _07699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08107_ _04503_ net1175 team_01_WB.instance_to_wrap.cpu.f0.state\[7\] _04577_ vssd1
+ vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__a31o_1
XFILLER_0_44_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09087_ net1011 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[13\] net930 vssd1
+ vssd1 vccd1 vccd1 _05427_ sky130_fd_sc_hd__and3_1
XANTENNA__12093__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08800__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08038_ net1665 net567 net345 team_01_WB.instance_to_wrap.cpu.f0.i\[17\] vssd1 vssd1
+ vccd1 vccd1 _03553_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_2_Left_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold850 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold861 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2396 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout596_X net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout975_A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11010__B net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1623_A team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold872 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[83\] vssd1 vssd1 vccd1 vccd1
+ net2407 sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[67\] vssd1 vssd1 vccd1 vccd1
+ net2418 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1303_X net1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold894 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[17\] vssd1 vssd1 vccd1 vccd1
+ net2429 sky130_fd_sc_hd__dlygate4sd3_1
X_10000_ _06339_ vssd1 vssd1 vccd1 vccd1 _06340_ sky130_fd_sc_hd__inv_2
X_09989_ _06325_ _06326_ _06327_ _06328_ vssd1 vssd1 vccd1 vccd1 _06329_ sky130_fd_sc_hd__or4_1
XANTENNA__10371__A1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1550 team_01_WB.instance_to_wrap.cpu.K0.code\[0\] vssd1 vssd1 vccd1 vccd1 net3085
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09513__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1561 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net3096 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_153_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11951_ net2161 net297 net478 vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__mux2_1
XANTENNA__09134__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout930_X net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1572 net149 vssd1 vssd1 vccd1 vccd1 net3107 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1583 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net3118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1594 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net3129 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_28_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10902_ _07003_ _07009_ net517 vssd1 vssd1 vccd1 vccd1 _07242_ sky130_fd_sc_hd__mux2_1
X_11882_ net3001 net280 net484 vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__mux2_1
X_14670_ net1224 vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_84_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08973__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11680__B net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10833_ _06220_ _07172_ vssd1 vssd1 vccd1 vccd1 _07173_ sky130_fd_sc_hd__or2_2
X_13621_ net186 _04059_ _04060_ net726 vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__a211o_1
XANTENNA__12268__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08619__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11623__A1 _07566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16340_ clknet_leaf_120_wb_clk_i net2758 _00323_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10764_ _05931_ net510 _06811_ net511 net542 net543 vssd1 vssd1 vccd1 vccd1 _07104_
+ sky130_fd_sc_hd__mux4_1
X_13552_ net196 net192 _07816_ _07861_ net643 vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_39_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12820__B1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10977__A3 _06526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12503_ net2667 net233 net407 vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__mux2_1
X_13483_ _03850_ _03851_ _03943_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__and3_1
X_16271_ clknet_leaf_159_wb_clk_i net1177 _00259_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.prev_BUSY_O
+ sky130_fd_sc_hd__dfrtp_1
X_10695_ _06902_ _07030_ _07032_ _07034_ _07026_ vssd1 vssd1 vccd1 vccd1 _07035_ sky130_fd_sc_hd__o41a_1
X_18010_ net637 vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11900__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15222_ net1258 vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__inv_2
X_12434_ net2168 net243 net417 vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__mux2_1
XANTENNA__13376__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15153_ net1419 vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__inv_2
X_12365_ net2705 net274 net425 vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11316_ team_01_WB.instance_to_wrap.cpu.f0.state\[8\] _07651_ vssd1 vssd1 vccd1 vccd1
+ _07653_ sky130_fd_sc_hd__or2_1
X_14104_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[53\] _04236_ _04244_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[101\]
+ _04390_ vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__a221o_1
X_15084_ net1259 vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12296_ net2436 net213 net431 vssd1 vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14035_ _04320_ _04321_ _04322_ _04324_ vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__or4_1
X_11247_ _06934_ _07524_ _07583_ vssd1 vssd1 vccd1 vccd1 _07587_ sky130_fd_sc_hd__a21oi_1
XANTENNA__15608__A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_55_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12731__S net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09752__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11178_ _07275_ _07515_ _07517_ _07514_ vssd1 vssd1 vccd1 vccd1 _07518_ sky130_fd_sc_hd__a211o_1
X_10129_ _06255_ _06410_ _06441_ _06468_ vssd1 vssd1 vccd1 vccd1 _06469_ sky130_fd_sc_hd__a211oi_4
X_15986_ net1363 vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__inv_2
X_17725_ clknet_leaf_156_wb_clk_i net873 _01666_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.state\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14937_ net1237 vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__inv_2
XANTENNA__09044__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17656_ clknet_leaf_4_wb_clk_i net1811 _01597_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11862__A1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14868_ net1379 vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16607_ clknet_leaf_41_wb_clk_i _02294_ _00590_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13819_ net2720 net832 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[12\]
+ sky130_fd_sc_hd__and2_1
X_17587_ clknet_leaf_124_wb_clk_i _03274_ _01546_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.code\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12178__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14799_ net1388 vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__inv_2
XANTENNA__13603__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11614__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16538_ clknet_leaf_6_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[4\]
+ _00521_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11090__A2 _05835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16469_ clknet_leaf_152_wb_clk_i _02223_ _00452_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11810__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09010_ net1095 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[9\] net914 vssd1
+ vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_94_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_103_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold102 net86 vssd1 vssd1 vccd1 vccd1 net1637 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 _01981_ vssd1 vssd1 vccd1 vccd1 net1648 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 _02013_ vssd1 vssd1 vccd1 vccd1 net1659 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09991__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold135 team_01_WB.instance_to_wrap.cpu.f0.write_data\[14\] vssd1 vssd1 vccd1 vccd1
+ net1670 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold146 team_01_WB.instance_to_wrap.cpu.f0.write_data\[26\] vssd1 vssd1 vccd1 vccd1
+ net1681 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 _02020_ vssd1 vssd1 vccd1 vccd1 net1692 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 _01997_ vssd1 vssd1 vccd1 vccd1 net1703 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold179 team_01_WB.instance_to_wrap.a1.ADR_I\[7\] vssd1 vssd1 vccd1 vccd1 net1714
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09912_ net556 _05264_ net377 vssd1 vssd1 vccd1 vccd1 _06252_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12641__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout604 _04151_ vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__clkbuf_4
Xfanout615 net616 vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__buf_4
Xfanout626 net627 vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09743__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout637 net179 vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__buf_2
X_09843_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[13\] net804 net784 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06183_ sky130_fd_sc_hd__a22o_1
Xfanout648 _04823_ vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08420__A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout659 _04813_ vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__buf_4
XANTENNA_fanout291_A _07941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout389_A _03569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09774_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[15\] net798 net785 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__a22o_1
XANTENNA__14095__A2 _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08725_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[5\] net672 _05045_ _05049_
+ _05051_ vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08849__A2 _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1298_A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08656_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[10\] net678 _04975_
+ _04977_ _04980_ vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_1_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09889__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08419__X _04759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12088__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08587_ net1031 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[15\] net909
+ vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__and3_1
XFILLER_0_152_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout723_A net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout344_X net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12802__B1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout511_X net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09208_ net1004 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[17\] net900
+ vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__and3_1
X_10480_ _06811_ _06813_ vssd1 vssd1 vccd1 vccd1 _06820_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09026__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09139_ net1110 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[14\] net913
+ vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08314__B net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12150_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[6\] net298 net454 vssd1
+ vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__mux2_1
XANTENNA__09982__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout880_X net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09129__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11101_ _07161_ _07440_ _07276_ vssd1 vssd1 vccd1 vccd1 _07441_ sky130_fd_sc_hd__a21o_1
X_12081_ net2005 net281 net460 vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__mux2_1
XANTENNA__12551__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold680 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2215 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold691 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2226 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08968__C net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13530__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11032_ _05417_ net341 vssd1 vssd1 vccd1 vccd1 _07372_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_34_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08330__A net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11541__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15840_ net1330 vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_139_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15771_ net1217 vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__inv_2
XANTENNA__13294__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12983_ net2337 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[111\] net856 vssd1 vssd1
+ vccd1 vccd1 _02142_ sky130_fd_sc_hd__mux2_1
X_17510_ clknet_leaf_83_wb_clk_i _03197_ _01493_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1380 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2915 sky130_fd_sc_hd__dlygate4sd3_1
X_14722_ net1189 vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__inv_2
Xhold1391 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2926 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11934_ net1973 net205 net475 vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17441_ clknet_leaf_54_wb_clk_i _03128_ _01424_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_14653_ net1270 vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__inv_2
X_11865_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[26\] net245 net485 vssd1
+ vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13597__A1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13604_ _03908_ _03900_ vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_107_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_107_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_17372_ clknet_leaf_58_wb_clk_i _03059_ _01355_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10816_ _05996_ net509 net508 net507 net549 net538 vssd1 vssd1 vccd1 vccd1 _07156_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_95_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11796_ net1975 net213 net491 vssd1 vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__mux2_1
X_14584_ net1354 vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__inv_2
XANTENNA__09265__A2 _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16323_ clknet_leaf_119_wb_clk_i _02077_ _00306_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13535_ net723 _07600_ net986 vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__a21oi_1
X_10747_ _06934_ _07065_ _07079_ _07086_ vssd1 vssd1 vccd1 vccd1 _07087_ sky130_fd_sc_hd__a211o_1
XFILLER_0_82_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11630__S net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16254_ clknet_leaf_141_wb_clk_i net1803 _00242_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10678_ _06963_ _06973_ _07016_ _06934_ _06997_ vssd1 vssd1 vccd1 vccd1 _07018_ sky130_fd_sc_hd__a221o_1
X_13466_ _05655_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] vssd1 vssd1
+ vccd1 vccd1 _03927_ sky130_fd_sc_hd__and2b_1
XANTENNA__16792__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14010__A2 _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10754__B net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15205_ net1275 vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__inv_2
X_12417_ net1792 net293 net421 vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__mux2_1
X_16185_ clknet_leaf_1_wb_clk_i _01945_ _00173_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13397_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] _05530_ vssd1 vssd1
+ vccd1 vccd1 _03858_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_58_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08776__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08776__B2 net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09973__B1 _06311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15136_ net1272 vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__inv_2
X_12348_ net2488 net302 net428 vssd1 vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15067_ net1254 vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__inv_2
XANTENNA__12461__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12279_ net2269 net227 net435 vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09725__B1 _06063_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14018_ _04295_ _04300_ _04305_ _04308_ vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_147_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09623__X _05963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15969_ net1403 vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__inv_2
XANTENNA__10099__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08510_ net1000 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[18\] net897 vssd1
+ vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__and3_1
XANTENNA__11805__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17708_ clknet_leaf_134_wb_clk_i _03392_ _01649_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_19_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09490_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[30\] net699 _05829_ net705
+ vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__a211o_1
XANTENNA__11835__A1 _07855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08700__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[7\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08441_ net1081 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[23\] net914
+ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__and3_1
X_17639_ clknet_leaf_0_wb_clk_i _03324_ _01580_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_33_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09502__C net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08372_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__nor2_2
XFILLER_0_73_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09110__D1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12636__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08415__A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14001__A2 _04226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10023__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09964__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12371__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13512__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout401 _03566_ vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__clkbuf_8
Xfanout412 _03563_ vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09716__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout423 net426 vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__clkbuf_8
Xfanout434 _07964_ vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__buf_4
XANTENNA_fanout673_A _04794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_6_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout445 _07959_ vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_92_Left_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout456 _07956_ vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09826_ net1143 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[13\] net965
+ vssd1 vssd1 vccd1 vccd1 _06166_ sky130_fd_sc_hd__and3_1
Xfanout467 net470 vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__buf_8
Xfanout478 _07950_ vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1001_X net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout489 _07947_ vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__buf_6
XANTENNA__12079__A1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10679__X _07019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13276__B1 _07650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09757_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[20\] net764 net623 vssd1
+ vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout840_A net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout461_X net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_5_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout559_X net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11715__S net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08708_ net1018 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[5\] net916 vssd1
+ vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__and3_1
X_09688_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[22\] net745 _06004_ _06008_
+ _06009_ vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__a2111o_1
X_08639_ net1020 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[10\] net902
+ vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__and3_1
XANTENNA__08309__B net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10558__C net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11650_ _07856_ _07857_ net611 vssd1 vssd1 vccd1 vccd1 _07858_ sky130_fd_sc_hd__mux2_4
XFILLER_0_49_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09247__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10601_ _06939_ _06940_ vssd1 vssd1 vccd1 vccd1 _06941_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11581_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] _07797_ vssd1 vssd1 vccd1
+ vccd1 _07798_ sky130_fd_sc_hd__and2_1
XANTENNA__12546__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10855__A net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13320_ net564 _07706_ _07731_ net828 vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__a31o_1
X_10532_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[31\] net654 net648 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06872_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13251_ _07686_ _07702_ vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__nor2_1
X_10463_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[26\] net798 net761 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06803_ sky130_fd_sc_hd__a22o_1
X_12202_ net2656 net271 net443 vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13182_ net1177 team_01_WB.instance_to_wrap.a1.prev_BUSY_O net835 vssd1 vssd1 vccd1
+ vccd1 _03738_ sky130_fd_sc_hd__and3b_2
XANTENNA__11211__C1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10394_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[16\] net821 _06732_ _06733_
+ vssd1 vssd1 vccd1 vccd1 _06734_ sky130_fd_sc_hd__a211o_1
XANTENNA_input67_A wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12133_ net1848 net205 net451 vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__mux2_1
XANTENNA__12281__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17990_ net635 vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_1
XANTENNA__13503__A1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09156__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12064_ net2516 net248 net461 vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__mux2_1
X_16941_ clknet_leaf_68_wb_clk_i _02628_ _00924_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11015_ _05594_ net508 vssd1 vssd1 vccd1 vccd1 _07355_ sky130_fd_sc_hd__xnor2_1
XANTENNA__16050__Q team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16872_ clknet_leaf_27_wb_clk_i _02559_ _00855_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout990 net995 vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__clkbuf_4
X_15823_ net1189 vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13267__B1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11625__S net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15754_ net1341 vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12966_ net1175 team_01_WB.instance_to_wrap.cpu.f0.state\[3\] vssd1 vssd1 vccd1 vccd1
+ _03718_ sky130_fd_sc_hd__nand2_1
XANTENNA__09486__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14705_ net1196 vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__inv_2
X_11917_ net2032 net279 net480 vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__mux2_1
X_15685_ net1289 vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__inv_2
X_12897_ net360 _03672_ net1036 vssd1 vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17424_ clknet_leaf_146_wb_clk_i _03111_ _01407_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14636_ net1388 vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__inv_2
X_11848_ net2497 net251 net490 vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__mux2_1
XANTENNA__09238__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17355_ clknet_leaf_11_wb_clk_i _03042_ _01338_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_14567_ net1406 vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11779_ net2393 net225 net495 vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11213__X _07553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16306_ clknet_leaf_100_wb_clk_i _02060_ _00289_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[29\]
+ sky130_fd_sc_hd__dfstp_1
X_13518_ net721 _07566_ net1074 vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__o21a_1
XANTENNA__12793__A2 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17286_ clknet_leaf_90_wb_clk_i _02973_ _01269_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14498_ net1363 vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__inv_2
X_16237_ clknet_leaf_133_wb_clk_i net1703 _00225_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__dfrtp_1
Xclkload11 clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload11/Y sky130_fd_sc_hd__inv_12
X_13449_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] _04946_ _03902_ vssd1
+ vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__a21o_1
Xclkload22 clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload22/Y sky130_fd_sc_hd__bufinv_16
Xclkload33 clknet_leaf_154_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload33/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_77_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_75_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xclkload44 clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload44/Y sky130_fd_sc_hd__inv_8
Xclkload55 clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload55/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__10005__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload66 clknet_leaf_65_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload66/Y sky130_fd_sc_hd__inv_6
XFILLER_0_23_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16168_ clknet_leaf_132_wb_clk_i net3093 _00156_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[31\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload77 clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload77/Y sky130_fd_sc_hd__inv_6
XANTENNA__10556__A1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09410__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload88 clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload88/Y sky130_fd_sc_hd__inv_6
XANTENNA__11596__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload99 clknet_leaf_131_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload99/Y sky130_fd_sc_hd__inv_6
X_15119_ net1388 vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_114_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12191__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08990_ net1087 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[8\] net926 vssd1
+ vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__and3_1
X_16099_ clknet_leaf_126_wb_clk_i _01874_ _00087_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10859__A2 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08921__A1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09611_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[24\] net789 net753 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__a22o_1
X_09542_ net1152 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[28\] net959
+ vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09477__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_924 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09473_ net1003 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[30\] net929 vssd1
+ vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout254_A net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08424_ net1082 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[23\] net935
+ vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08355_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[30\] net817 net759 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[30\]
+ _04694_ vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12366__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13861__A_N net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13430__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout421_A net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10244__B1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout519_A net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12784__A2 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload5 clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload5/Y sky130_fd_sc_hd__inv_4
X_08286_ net1170 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__or3b_4
XFILLER_0_33_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10795__A1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1330_A net1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1428_A net1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13733__A1 team_01_WB.instance_to_wrap.cpu.DM0.dhit vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13733__B2 team_01_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08432__X _04772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout790_A _04654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09401__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout888_A _04799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11744__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1536_A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08151__Y _04621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1207 net1304 vssd1 vssd1 vccd1 vccd1 net1207 sky130_fd_sc_hd__buf_2
XANTENNA__13497__B1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12889__X _03667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout220 _07831_ vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__buf_2
Xfanout1218 net1219 vssd1 vssd1 vccd1 vccd1 net1218 sky130_fd_sc_hd__buf_4
Xfanout1229 net1304 vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__clkbuf_4
Xfanout231 net232 vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__buf_2
XANTENNA_fanout676_X net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout242 net243 vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__buf_2
Xfanout253 net256 vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__buf_2
Xfanout264 _07880_ vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout275 _07851_ vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__clkbuf_2
Xfanout286 _07896_ vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__clkbuf_2
Xfanout297 _07921_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__clkbuf_2
X_09809_ _06141_ _06142_ _06143_ _06148_ vssd1 vssd1 vccd1 vccd1 _06149_ sky130_fd_sc_hd__or4_1
XANTENNA__09704__A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout843_X net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12820_ net364 _03641_ _03642_ net1062 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__a32o_1
X_12751_ net1040 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[25\] vssd1 vssd1 vccd1
+ vccd1 _03595_ sky130_fd_sc_hd__or2_2
XFILLER_0_57_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11702_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] _07803_ vssd1 vssd1
+ vccd1 vccd1 _07899_ sky130_fd_sc_hd__or2_1
X_15470_ net1298 vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__inv_2
X_12682_ net2329 net312 net390 vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08981__C net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14421_ net1335 vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11633_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[25\] net715 net615 vssd1 vssd1
+ vccd1 vccd1 _07844_ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12276__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17140_ clknet_leaf_21_wb_clk_i _02827_ _01123_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_14352_ net1326 vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11564_ team_01_WB.instance_to_wrap.cpu.K0.count\[1\] team_01_WB.instance_to_wrap.cpu.K0.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__nand2_1
XANTENNA__10786__A1 _04919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13303_ team_01_WB.instance_to_wrap.cpu.f0.i\[20\] net610 _07707_ team_01_WB.instance_to_wrap.cpu.f0.i\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__a31o_1
X_17071_ clknet_leaf_35_wb_clk_i _02758_ _01054_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10515_ _06847_ _06848_ _06853_ _06854_ vssd1 vssd1 vccd1 vccd1 _06855_ sky130_fd_sc_hd__or4_2
XFILLER_0_150_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14283_ net1336 vssd1 vssd1 vccd1 vccd1 _00077_ sky130_fd_sc_hd__inv_2
X_11495_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[15\] net580 vssd1 vssd1 vccd1
+ vccd1 _07775_ sky130_fd_sc_hd__nand2_1
XANTENNA__09928__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16022_ net1340 vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13234_ net2871 net352 net348 team_01_WB.instance_to_wrap.cpu.f0.i\[16\] vssd1 vssd1
+ vccd1 vccd1 _01916_ sky130_fd_sc_hd__a22o_1
X_10446_ net1147 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[26\] net974
+ vssd1 vssd1 vccd1 vccd1 _06786_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_94_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10538__A1 net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10377_ net1143 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[16\] net966
+ vssd1 vssd1 vccd1 vccd1 _06717_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13165_ net110 net849 net841 net1798 vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_72_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12116_ net2760 net277 net455 vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__mux2_1
X_13096_ net50 net39 net64 net61 vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__or4_1
X_17973_ net1488 vssd1 vssd1 vccd1 vccd1 la_data_out[15] sky130_fd_sc_hd__buf_2
XANTENNA__13488__B1 _05780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12799__X _03628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_144_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12047_ net1767 net249 net466 vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__mux2_1
X_16924_ clknet_leaf_59_wb_clk_i _02611_ _00907_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_140_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16855_ clknet_leaf_17_wb_clk_i _02542_ _00838_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_140_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15806_ net1206 vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_122_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_122_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_148_Left_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16786_ clknet_leaf_145_wb_clk_i _02473_ _00769_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13998_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[3\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\]
+ _04237_ vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__and3b_1
X_15737_ net1238 vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__inv_2
XANTENNA__09052__C net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11266__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12949_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[7\] net1041 vssd1 vssd1 vccd1
+ vccd1 _03709_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10198__C net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15668_ net1379 vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08891__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17407_ clknet_leaf_39_wb_clk_i _03094_ _01390_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14619_ net1342 vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__inv_2
XANTENNA__12186__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15599_ net1388 vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08140_ _04606_ _04607_ _04608_ _04609_ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__or4_1
XFILLER_0_16_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17338_ clknet_leaf_78_wb_clk_i _03025_ _01321_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17486__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10777__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload100 clknet_leaf_132_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload100/Y sky130_fd_sc_hd__inv_6
X_08071_ _04515_ _04523_ _04537_ _04546_ vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__or4_1
XFILLER_0_114_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload111 clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload111/Y sky130_fd_sc_hd__inv_6
X_17269_ clknet_leaf_111_wb_clk_i _02956_ _01252_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload122 clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload122/Y sky130_fd_sc_hd__clkinv_2
Xclkload133 clknet_leaf_92_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload133/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__09495__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload144 clknet_leaf_85_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload144/Y sky130_fd_sc_hd__inv_6
XANTENNA__09919__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13191__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08412__B net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08973_ net1007 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[8\] net926 vssd1
+ vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__and3_1
Xhold17 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[5\] vssd1 vssd1 vccd1 vccd1
+ net1552 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[17\] vssd1 vssd1 vccd1 vccd1 net1563
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 _02026_ vssd1 vssd1 vccd1 vccd1 net1574 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1009_A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout371_A _06738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout469_A net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11065__A2_N net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09525_ _05855_ _05860_ _05864_ vssd1 vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__nor3_1
XFILLER_0_78_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout636_A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1378_A net1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_5_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09456_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[29\] net697 net691 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[29\]
+ _05786_ vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09870__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08407_ _04738_ _04745_ vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__and2b_1
XFILLER_0_47_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12096__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout803_A _04643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout424_X net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09387_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] net710 _04841_ vssd1 vssd1
+ vccd1 vccd1 _05727_ sky130_fd_sc_hd__a21o_1
XANTENNA__13403__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10217__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08338_ net1139 net965 vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__and2_4
XFILLER_0_85_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09622__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07985__Y _04483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08269_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[12\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[4\]
+ net1045 vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10300_ net505 _06638_ vssd1 vssd1 vccd1 vccd1 _06640_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11280_ _07054_ _07497_ _07614_ _06963_ _07619_ vssd1 vssd1 vccd1 vccd1 _07620_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout793_X net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10231_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[9\] net744 net741 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06571_ sky130_fd_sc_hd__a22o_1
X_10162_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] net626 vssd1 vssd1 vccd1
+ vccd1 _06502_ sky130_fd_sc_hd__nand2_1
XANTENNA__09137__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1004 net1015 vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__buf_2
Xfanout1015 _04490_ vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__clkbuf_2
Xfanout1026 net1030 vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__buf_2
X_10093_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[7\] net814 net779 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[7\]
+ _06411_ vssd1 vssd1 vccd1 vccd1 _06433_ sky130_fd_sc_hd__a221o_1
Xfanout1037 net1041 vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__clkbuf_4
X_14970_ net1314 vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__inv_2
Xfanout1048 net1049 vssd1 vssd1 vccd1 vccd1 net1048 sky130_fd_sc_hd__clkbuf_4
Xfanout1059 team_01_WB.instance_to_wrap.cpu.SR1.enable vssd1 vssd1 vccd1 vccd1 net1059
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_156_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08976__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13921_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[13\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[12\]
+ _04212_ vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__and3_1
XFILLER_0_156_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16640_ clknet_leaf_46_wb_clk_i _02327_ _00623_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08361__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13852_ net1179 net1066 net1708 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[13\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_92_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12803_ net1762 net640 net608 _03630_ vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_48_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16571_ clknet_leaf_68_wb_clk_i _02258_ _00554_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_13783_ _04162_ _01835_ _04166_ _04159_ vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__o211a_1
XANTENNA__10867__X _07207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10995_ net563 net337 _07334_ vssd1 vssd1 vccd1 vccd1 _07335_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11903__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15522_ net1351 vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__inv_2
X_12734_ net1953 net638 _03582_ net606 vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09861__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15453_ net1240 vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__inv_2
X_12665_ net2547 net242 net389 vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12748__A2 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14404_ net1360 vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11616_ net615 _07830_ _07829_ vssd1 vssd1 vccd1 vccd1 _07831_ sky130_fd_sc_hd__o21ai_4
XANTENNA__11405__C1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15384_ net1214 vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_96_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09613__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12596_ net2226 net273 net397 vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11698__X _07896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17123_ clknet_leaf_25_wb_clk_i _02810_ _01106_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14335_ net1341 vssd1 vssd1 vccd1 vccd1 _00129_ sky130_fd_sc_hd__inv_2
X_11547_ net1995 net1174 vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_133_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17054_ clknet_leaf_80_wb_clk_i _02741_ _01037_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold509 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2044 sky130_fd_sc_hd__dlygate4sd3_1
X_14266_ net1224 vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__inv_2
X_11478_ net367 _07766_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[24\] net875
+ vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_111_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16005_ net1328 vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_111_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13217_ net566 _03740_ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__or2_1
X_10429_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[27\] net782 _06755_ _06759_
+ _06762_ vssd1 vssd1 vccd1 vccd1 _06769_ sky130_fd_sc_hd__a2111o_1
X_14197_ net1588 _04462_ net1428 vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13148_ net1616 net846 net839 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[28\] vssd1
+ vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__a22o_1
XANTENNA__09047__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17956_ net1471 vssd1 vssd1 vccd1 vccd1 irq[1] sky130_fd_sc_hd__buf_2
XANTENNA__14250__A net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13079_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[7\] net2883 net858 vssd1 vssd1
+ vccd1 vccd1 _02046_ sky130_fd_sc_hd__mux2_1
Xhold1209 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2744 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08886__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09344__A net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16907_ clknet_leaf_10_wb_clk_i _02594_ _00890_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_17887_ net107 vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_109_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08352__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16838_ clknet_leaf_73_wb_clk_i _02525_ _00821_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_68_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12436__A1 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16769_ clknet_leaf_57_wb_clk_i _02456_ _00752_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11813__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09310_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[22\] net664 _05627_
+ _05629_ _05641_ vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_76_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09241_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[21\] net671 net648 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09510__C net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_90_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_118_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09172_ net1010 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[16\] net910
+ vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12739__A2 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08123_ _04480_ team_01_WB.instance_to_wrap.cpu.f0.num\[14\] team_01_WB.instance_to_wrap.cpu.f0.num\[13\]
+ _04481_ vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_16_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12644__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08812__B1 _05116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout217_A _07835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08054_ team_01_WB.instance_to_wrap.cpu.K0.code\[7\] team_01_WB.instance_to_wrap.cpu.K0.code\[6\]
+ team_01_WB.instance_to_wrap.cpu.K0.code\[4\] team_01_WB.instance_to_wrap.cpu.K0.code\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__or4b_2
XANTENNA__13164__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11175__A1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1126_A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10367__A1_N net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout586_A net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08591__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08956_ _05292_ _05293_ _05294_ _05295_ vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__or4_1
XANTENNA__08796__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08879__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout753_A net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08887_ net1107 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[2\] net924 vssd1
+ vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout374_X net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10150__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout920_A net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10438__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09508_ net1149 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[29\] net979
+ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__and3_1
X_10780_ net515 _07105_ vssd1 vssd1 vccd1 vccd1 _07120_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09843__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09439_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[28\] net703 _05774_ _05778_
+ vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__o22a_2
XANTENNA_fanout806_X net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08317__B net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12450_ net2853 net294 net417 vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__mux2_1
X_11401_ _07696_ _07714_ team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1 vccd1
+ vccd1 _07724_ sky130_fd_sc_hd__a21o_1
XFILLER_0_90_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12381_ net1932 net302 net424 vssd1 vssd1 vccd1 vccd1 _02615_ sky130_fd_sc_hd__mux2_1
XANTENNA__12554__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08604__Y _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14120_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[86\] _04251_ _04255_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[118\]
+ _04397_ vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__a221o_1
X_11332_ _07664_ net2086 _07655_ vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08333__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10582__B _06920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14054__B _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13155__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14051_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[75\] _04235_ _04250_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[123\]
+ _04339_ vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__a221o_1
X_11263_ net528 _07106_ vssd1 vssd1 vccd1 vccd1 _07603_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_45_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_120_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13002_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[84\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[92\]
+ net855 vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__mux2_1
X_10214_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[8\] net748 _06537_ _06541_
+ _06543_ vssd1 vssd1 vccd1 vccd1 _06554_ sky130_fd_sc_hd__a2111o_1
X_11194_ _07058_ _07080_ net515 vssd1 vssd1 vccd1 vccd1 _07534_ sky130_fd_sc_hd__mux2_1
X_17810_ clknet_leaf_123_wb_clk_i net3087 _01750_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[80\]
+ sky130_fd_sc_hd__dfrtp_1
X_10145_ _06481_ _06482_ _06483_ _06484_ vssd1 vssd1 vccd1 vccd1 _06485_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_37_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09164__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17741_ clknet_leaf_96_wb_clk_i _03417_ _01681_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10076_ net1138 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[7\] net965 vssd1
+ vssd1 vccd1 vccd1 _06416_ sky130_fd_sc_hd__and3_1
X_14953_ net1288 vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_89_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13904_ _04204_ net571 _04203_ vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__and3b_1
X_17672_ clknet_leaf_0_wb_clk_i _03357_ _01613_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10103__A net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14884_ net1217 vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__inv_2
XANTENNA__10141__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16623_ clknet_leaf_36_wb_clk_i _02310_ _00606_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13835_ net1668 net830 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[28\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_134_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13414__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16554_ clknet_leaf_0_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[20\]
+ _00537_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13766_ _04154_ vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__inv_2
XANTENNA__13091__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10978_ _06438_ net372 net551 vssd1 vssd1 vccd1 vccd1 _07318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08508__A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09834__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15505_ net1393 vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__inv_2
X_12717_ net2340 net318 net386 vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16485_ clknet_leaf_141_wb_clk_i _02239_ _00468_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_135_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13697_ _04110_ _04111_ _04119_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[15\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_150_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15436_ net1260 vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12648_ net2721 net295 net393 vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_84_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_5_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_152_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15367_ net1391 vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__inv_2
XANTENNA__12464__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12579_ net2021 net300 net400 vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17106_ clknet_leaf_145_wb_clk_i _02793_ _01089_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_14318_ net1327 vssd1 vssd1 vccd1 vccd1 _00112_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08270__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold306 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[28\] vssd1 vssd1 vccd1 vccd1
+ net1841 sky130_fd_sc_hd__dlygate4sd3_1
X_15298_ net1318 vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__inv_2
Xhold317 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1852 sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1863 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13146__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold339 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[3\] vssd1 vssd1 vccd1 vccd1 net1874
+ sky130_fd_sc_hd__dlygate4sd3_1
X_17037_ clknet_leaf_109_wb_clk_i _02724_ _01020_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_14249_ net1218 vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__inv_2
Xfanout808 net810 vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout819 _04632_ vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__buf_6
X_08810_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[0\] net702 _05133_ _05149_
+ vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__o22a_4
XANTENNA__11808__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09790_ net376 net342 _05492_ net560 vssd1 vssd1 vccd1 vccd1 _06130_ sky130_fd_sc_hd__a31o_1
XANTENNA__10380__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1006 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[43\] vssd1 vssd1 vccd1 vccd1
+ net2541 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1017 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2552 sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ net1099 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[4\] net916 vssd1
+ vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__and3_1
X_17939_ net1454 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
XFILLER_0_139_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1028 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2563 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17674__CLK clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12657__A1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1039 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2574 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09505__C net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1390 net1391 vssd1 vssd1 vccd1 vccd1 net1390 sky130_fd_sc_hd__buf_4
X_08672_ net1085 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[7\] net939 vssd1
+ vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08730__C1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12639__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08418__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10667__B _06250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10840__A0 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09224_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[17\] net702 _05561_ _05563_
+ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__o22a_4
XFILLER_0_57_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14031__B1 _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09155_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[16\] net620 net593 vssd1 vssd1
+ vccd1 vccd1 _05495_ sky130_fd_sc_hd__a21o_1
XANTENNA__12374__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout501_A net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1243_A net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08106_ _04511_ _04575_ _04576_ net1041 vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__o31a_1
X_09086_ net1011 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[13\] _04779_
+ vssd1 vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08037_ net1646 net567 net345 team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1
+ vccd1 vccd1 _03554_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1031_X net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold840 team_01_WB.instance_to_wrap.cpu.c0.count\[2\] vssd1 vssd1 vccd1 vccd1 net2375
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11148__A1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17974__1489 vssd1 vssd1 vccd1 vccd1 _17974__1489/HI net1489 sky130_fd_sc_hd__conb_1
Xhold851 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2386 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1129_X net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13542__C1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold862 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2397 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07992__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold873 _03489_ vssd1 vssd1 vccd1 vccd1 net2408 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold884 _03473_ vssd1 vssd1 vccd1 vccd1 net2419 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08440__X _04780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout870_A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout491_X net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold895 _03431_ vssd1 vssd1 vccd1 vccd1 net2430 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11718__S net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout968_A _04648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08564__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09988_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[2\] net796 net789 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06328_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_129_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08939_ net1027 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[6\] net881 vssd1
+ vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__and3_1
XANTENNA__12648__A1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_150_Right_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout756_X net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10659__A0 _06158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1540 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 net3075
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1551 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[72\] vssd1 vssd1 vccd1 vccd1
+ net3086 sky130_fd_sc_hd__dlygate4sd3_1
X_11950_ net2483 net278 net476 vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__mux2_1
Xhold1562 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net3097 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10123__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1573 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net3108 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_28_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1584 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net3119 sky130_fd_sc_hd__dlygate4sd3_1
X_10901_ net523 _07240_ vssd1 vssd1 vccd1 vccd1 _07241_ sky130_fd_sc_hd__or2_1
Xhold1595 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net3130 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11881_ net2663 net249 net486 vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout923_X net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12549__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17702__Q team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13620_ net197 net193 _07804_ _07903_ net643 vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__o2111a_1
X_10832_ _06469_ _06472_ _06597_ _06603_ vssd1 vssd1 vccd1 vccd1 _07172_ sky130_fd_sc_hd__o31a_1
XFILLER_0_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08328__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13551_ _03932_ _04001_ vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__xnor2_1
X_10763_ _06958_ _07099_ _07102_ _07098_ vssd1 vssd1 vccd1 vccd1 _07103_ sky130_fd_sc_hd__a211o_1
XANTENNA__12820__A1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12502_ net2555 net237 net407 vssd1 vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10831__B1 _07170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16270_ clknet_leaf_124_wb_clk_i _02030_ _00258_ vssd1 vssd1 vccd1 vccd1 team_01_WB.EN_VAL_REG
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_137_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14022__B1 _04241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13482_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] _05679_ _05705_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\]
+ _03941_ vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__a221o_1
X_10694_ _06906_ _07033_ vssd1 vssd1 vccd1 vccd1 _07034_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15221_ net1282 vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__inv_2
X_12433_ net2550 net202 net415 vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12284__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15152_ net1273 vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12364_ net1785 net209 net425 vssd1 vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16053__Q team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14103_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[45\] _04246_ _04251_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[85\]
+ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13128__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11315_ team_01_WB.instance_to_wrap.cpu.f0.state\[8\] _07651_ vssd1 vssd1 vccd1 vccd1
+ _07652_ sky130_fd_sc_hd__nor2_2
X_15083_ net1423 vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_112_Left_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12295_ net1908 net214 net431 vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14034_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[26\] _04243_ _04254_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[98\]
+ _04323_ vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__a221o_1
X_11246_ net556 _07528_ _07582_ _07345_ _07585_ vssd1 vssd1 vccd1 vccd1 _07586_ sky130_fd_sc_hd__o221a_1
XFILLER_0_129_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08555__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13409__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11177_ net531 _07445_ _07516_ net328 vssd1 vssd1 vccd1 vccd1 _07517_ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10362__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10128_ net372 _06467_ vssd1 vssd1 vccd1 vccd1 _06468_ sky130_fd_sc_hd__and2_1
X_15985_ net1410 vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17724_ clknet_leaf_156_wb_clk_i _00006_ _01665_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.state\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_14936_ net1210 vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__inv_2
X_10059_ net552 _06398_ vssd1 vssd1 vccd1 vccd1 _06399_ sky130_fd_sc_hd__or2_2
XANTENNA__10114__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_121_Left_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14867_ net1404 vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__inv_2
X_17655_ clknet_leaf_5_wb_clk_i net1721 _01596_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12459__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16606_ clknet_leaf_80_wb_clk_i _02293_ _00589_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13818_ net2150 net833 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[11\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_102_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17586_ clknet_leaf_130_wb_clk_i _03273_ _01545_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.code\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09268__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14798_ net1291 vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__inv_2
XANTENNA__09807__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16537_ clknet_leaf_6_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[3\]
+ _00520_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_154_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09060__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11614__A2 _07056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13749_ _04115_ team_01_WB.instance_to_wrap.cpu.c0.next_count\[16\] _04138_ team_01_WB.instance_to_wrap.cpu.c0.next_count\[0\]
+ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_atmax sky130_fd_sc_hd__and4b_1
XANTENNA__12811__A1 _07323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16468_ clknet_leaf_14_wb_clk_i _02222_ _00451_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14013__B1 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11599__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15419_ net1252 vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__inv_2
XANTENNA__12194__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16399_ clknet_leaf_91_wb_clk_i net1743 _00382_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_130_Left_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold103 _01999_ vssd1 vssd1 vccd1 vccd1 net1638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[121\] vssd1 vssd1 vccd1 vccd1
+ net1649 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13119__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold125 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 net1660
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12922__S net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold136 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[14\] vssd1 vssd1 vccd1 vccd1
+ net1671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 team_01_WB.instance_to_wrap.cpu.c0.count\[0\] vssd1 vssd1 vccd1 vccd1 net1682
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 net129 vssd1 vssd1 vccd1 vccd1 net1693 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ _06250_ vssd1 vssd1 vccd1 vccd1 _06251_ sky130_fd_sc_hd__inv_2
Xhold169 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net1704 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12878__A1 _03659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout605 _04151_ vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__clkbuf_2
Xfanout616 _07635_ vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09842_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[13\] net786 net741 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[13\]
+ _06181_ vssd1 vssd1 vccd1 vccd1 _06182_ sky130_fd_sc_hd__a221o_1
XANTENNA__09075__Y _05415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout627 _04627_ vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__clkbuf_8
Xfanout638 _03572_ vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__buf_2
Xfanout649 _04823_ vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08420__B net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10353__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[15\] net792 net751 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[15\]
+ _06112_ vssd1 vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout284_A _07896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08724_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[5\] net700 net667 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__a22o_1
XANTENNA__10105__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09532__A net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08655_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[10\] net669 _04989_ _04993_
+ _04994_ vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_1_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout451_A _07957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12369__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout549_A _05151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09259__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08586_ net1031 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[15\] net942 vssd1
+ vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12802__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout337_X net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout716_A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07987__A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1079_X net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14004__B1 _04266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09207_ net1082 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[17\] net904
+ vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout504_X net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09138_ net1110 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[14\] net908
+ vssd1 vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__and3_1
XANTENNA__09431__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07993__Y _04491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09069_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[12\] net691 _05384_ _05395_
+ _05403_ vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_102_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11100_ _06921_ _07160_ vssd1 vssd1 vccd1 vccd1 _07440_ sky130_fd_sc_hd__or2_1
XANTENNA__09707__A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12080_ net2428 net249 net462 vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__mux2_1
XANTENNA__12869__A1 _06881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold670 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[25\] vssd1 vssd1 vccd1 vccd1
+ net2205 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout873_X net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold681 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2216 sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2227 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13530__A2 _07579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11031_ _07369_ _07370_ vssd1 vssd1 vccd1 vccd1 _07371_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_34_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11541__B2 net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15770_ net1217 vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_51_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13294__A1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12982_ net2710 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[112\] net853 vssd1 vssd1
+ vccd1 vccd1 _02143_ sky130_fd_sc_hd__mux2_1
Xhold1370 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2905 sky130_fd_sc_hd__dlygate4sd3_1
X_14721_ net1188 vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__inv_2
XANTENNA_input12_A DAT_I[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1381 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2916 sky130_fd_sc_hd__dlygate4sd3_1
X_11933_ net2554 net274 net477 vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__mux2_1
Xhold1392 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2927 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12279__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17440_ clknet_leaf_45_wb_clk_i _03127_ _01423_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14652_ net1314 vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__inv_2
X_11864_ net1960 net213 net483 vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13603_ net987 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] _04044_ _04045_
+ vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__a22o_1
X_17371_ clknet_leaf_74_wb_clk_i _03058_ _01354_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10815_ _06106_ _06744_ _06747_ vssd1 vssd1 vccd1 vccd1 _07155_ sky130_fd_sc_hd__nand3_1
XANTENNA__13597__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16048__Q team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14583_ net1402 vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__inv_2
X_11795_ net2035 net217 net493 vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__mux2_1
XANTENNA__11911__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16322_ clknet_leaf_101_wb_clk_i _02076_ _00305_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[45\]
+ sky130_fd_sc_hd__dfstp_1
X_13534_ net186 _03986_ _03987_ net723 vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__a211o_1
X_10746_ net523 _07082_ _07083_ _05263_ _07085_ vssd1 vssd1 vccd1 vccd1 _07086_ sky130_fd_sc_hd__o221a_1
XFILLER_0_125_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16253_ clknet_leaf_152_wb_clk_i net1659 _00241_ vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_147_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_147_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_82_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13465_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] _04842_ vssd1 vssd1
+ vccd1 vccd1 _03926_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10677_ net556 _06858_ _06921_ vssd1 vssd1 vccd1 vccd1 _07017_ sky130_fd_sc_hd__a21oi_4
XANTENNA__11212__A _07550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15204_ net1218 vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12416_ net2766 net299 net422 vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16184_ clknet_leaf_6_wb_clk_i _01944_ _00172_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13396_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] _05530_ vssd1 vssd1
+ vccd1 vccd1 _03857_ sky130_fd_sc_hd__and2_1
XANTENNA__09422__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09973__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15135_ net1318 vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__inv_2
X_12347_ net2989 net281 net428 vssd1 vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13506__C1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15066_ net1370 vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__inv_2
X_12278_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[12\] net287 net437 vssd1
+ vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14017_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[49\] _04236_ _04290_ _04307_
+ _04152_ vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09725__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11229_ _05965_ _07568_ _05934_ vssd1 vssd1 vccd1 vccd1 _07569_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_147_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11532__B2 net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09055__C net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13285__A1 _04621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09489__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15968_ net1354 vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__inv_2
XANTENNA__08894__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17707_ clknet_leaf_134_wb_clk_i _03391_ _01648_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[28\]
+ sky130_fd_sc_hd__dfrtp_4
X_14919_ net1390 vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__inv_2
XANTENNA__12189__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08697__D1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10498__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15899_ net1367 vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_121_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08700__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08440_ net1097 net916 vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__and2_1
X_17638_ clknet_leaf_0_wb_clk_i _03323_ _01579_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17973__1488 vssd1 vssd1 vccd1 vccd1 _17973__1488/HI net1488 sky130_fd_sc_hd__conb_1
X_08371_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[3\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[2\]
+ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[1\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_92_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17569_ clknet_leaf_87_wb_clk_i _03256_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11821__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12796__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire886_A _04803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09413__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_3_0_wb_clk_i_X clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08767__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12652__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11771__A1 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1039_A net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout402 _03566_ vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout499_A net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout413 _03563_ vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__buf_6
XANTENNA__10025__X _06365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout424 net426 vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1206_A net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout435 net438 vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__buf_6
Xfanout446 _07959_ vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__buf_4
XANTENNA__11523__B2 team_01_WB.instance_to_wrap.cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12720__B1 net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09825_ _06134_ _06164_ vssd1 vssd1 vccd1 vccd1 _06165_ sky130_fd_sc_hd__or2_1
XANTENNA_input4_A DAT_I[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout457 _07956_ vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__clkbuf_8
Xfanout468 net470 vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout666_A _04804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout479 _07949_ vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__buf_6
X_09756_ net768 _06089_ _06093_ _06095_ vssd1 vssd1 vccd1 vccd1 _06096_ sky130_fd_sc_hd__nor4_1
XANTENNA__13276__A1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08707_ net1018 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[5\] net919 vssd1
+ vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__and3_1
X_09687_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[22\] net782 net759 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__a22o_1
XANTENNA__12099__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout454_X net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout833_A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08638_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[10\] net908
+ vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11016__B net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08569_ net999 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[19\] net878 vssd1
+ vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout719_X net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12787__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10600_ net546 net339 vssd1 vssd1 vccd1 vccd1 _06940_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11580_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\]
+ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1 vccd1 vccd1 _07797_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_107_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10855__B net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10531_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[31\] net693 net686 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06871_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13250_ net2511 net353 net349 team_01_WB.instance_to_wrap.cpu.f0.i\[0\] vssd1 vssd1
+ vccd1 vccd1 _01900_ sky130_fd_sc_hd__a22o_1
X_10462_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[26\] net792 net773 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06802_ sky130_fd_sc_hd__a22o_1
XANTENNA__09404__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout990_X net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12201_ net2042 net241 net445 vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__mux2_1
X_13181_ team_01_WB.instance_to_wrap.a1.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1
+ _03737_ sky130_fd_sc_hd__nand2_1
XANTENNA__12562__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10393_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[16\] net803 net754 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06733_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11762__A1 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12132_ net2325 net274 net453 vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08341__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10970__C1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16940_ clknet_leaf_16_wb_clk_i _02627_ _00923_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_12063_ net2003 net212 net459 vssd1 vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11514__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10317__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11014_ _05595_ net508 vssd1 vssd1 vccd1 vccd1 _07354_ sky130_fd_sc_hd__nand2_1
X_16871_ clknet_leaf_106_wb_clk_i _02558_ _00854_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15174__A net1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout980 _04633_ vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__buf_4
XANTENNA__11906__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout991 net992 vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__clkbuf_2
X_15822_ net1190 vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_142_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09172__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15753_ net1341 vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__inv_2
X_12965_ net1770 net871 net358 _03717_ vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__a22o_1
XANTENNA__09603__C net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11916_ net2422 net302 net480 vssd1 vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__mux2_1
XANTENNA__15902__A net1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14704_ net1196 vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__inv_2
X_15684_ net1219 vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__inv_2
X_12896_ _04837_ net577 vssd1 vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14635_ net1291 vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__inv_2
X_17423_ clknet_leaf_33_wb_clk_i _03110_ _01406_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11847_ net2545 net225 net487 vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12778__B1 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17354_ clknet_leaf_10_wb_clk_i _03041_ _01337_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_14566_ net1401 vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__inv_2
X_11778_ net2310 net284 net497 vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08516__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13517_ net187 _03972_ _03973_ net727 vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__a211o_1
X_16305_ clknet_leaf_118_wb_clk_i _02059_ _00288_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[28\]
+ sky130_fd_sc_hd__dfstp_1
X_17285_ clknet_leaf_49_wb_clk_i _02972_ _01268_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10729_ _06920_ _06928_ vssd1 vssd1 vccd1 vccd1 _07069_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13990__A2 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14497_ net1364 vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16236_ clknet_leaf_133_wb_clk_i net1795 _00224_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__dfrtp_1
Xclkload12 clknet_leaf_155_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload12/Y sky130_fd_sc_hd__clkinv_16
X_13448_ _03904_ _03907_ _03908_ vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__nand3_1
Xclkload23 clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload23/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_77_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload34 clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload34/Y sky130_fd_sc_hd__inv_6
Xclkload45 clknet_leaf_35_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload45/Y sky130_fd_sc_hd__inv_6
Xclkload56 clknet_leaf_47_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload56/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__12472__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16167_ clknet_leaf_131_wb_clk_i _01930_ _00155_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13379_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] _05834_ vssd1 vssd1
+ vccd1 vccd1 _03840_ sky130_fd_sc_hd__and2b_1
XANTENNA__14253__A net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload67 clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload67/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_149_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload78 clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload78/Y sky130_fd_sc_hd__inv_6
XFILLER_0_51_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08889__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15118_ net1298 vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_114_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload89 clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload89/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_114_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16098_ clknet_leaf_126_wb_clk_i _01873_ _00086_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_15049_ net1287 vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_44_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09174__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10859__A3 _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11816__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09610_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[24\] net757 _05936_ _05942_
+ _05945_ vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08921__A2 _05258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09541_ net997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[28\] _04640_
+ vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09472_ net1080 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[30\] net901
+ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__and3_1
XFILLER_0_149_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08423_ net1108 net936 vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__and2_1
XANTENNA__12647__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12769__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout247_A _07842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08354_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[30\] net786 net734 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__a22o_1
XANTENNA__13430__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08426__A net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload6 clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload6/Y sky130_fd_sc_hd__inv_6
X_08285_ _04623_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[3\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__or3b_1
XANTENNA__13981__A2 _04265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout414_A _03563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1156_A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13194__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12382__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10691__A _05190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout202_X net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14163__A net1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08799__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout783_A net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13497__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1208 net1209 vssd1 vssd1 vccd1 vccd1 net1208 sky130_fd_sc_hd__buf_4
Xfanout210 net211 vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__buf_2
XFILLER_0_10_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1219 net1223 vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__buf_2
Xfanout221 net224 vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1209_X net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout232 _07884_ vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09165__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout243 net244 vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__buf_2
XFILLER_0_100_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout254 net256 vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__buf_2
Xfanout265 net266 vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout669_X net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout276 net279 vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__buf_2
XANTENNA__08912__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout287 _07896_ vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__buf_1
X_09808_ _06144_ _06145_ _06146_ _06147_ vssd1 vssd1 vccd1 vccd1 _06148_ sky130_fd_sc_hd__or4_1
Xfanout298 _07921_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__buf_2
XANTENNA__10180__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_15__f_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_15__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__13249__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_119_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09739_ net1145 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[20\] net970
+ vssd1 vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__and3_1
X_12750_ net1034 _07579_ vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11701_ net718 _07207_ net615 _07897_ vssd1 vssd1 vccd1 vccd1 _07898_ sky130_fd_sc_hd__o211a_1
X_12681_ net2314 net292 net389 vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__mux2_1
XANTENNA__12557__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14420_ net1307 vssd1 vssd1 vccd1 vccd1 _00214_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11632_ net715 _07579_ vssd1 vssd1 vccd1 vccd1 _07843_ sky130_fd_sc_hd__nand2_1
XANTENNA__08336__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08979__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14351_ net1338 vssd1 vssd1 vccd1 vccd1 _00145_ sky130_fd_sc_hd__inv_2
XANTENNA__11432__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_53_926 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11563_ net3083 net1182 net34 vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__a21o_1
XANTENNA__10786__A2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13302_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[24\] net825 _03783_ _03785_
+ vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__o22a_1
XFILLER_0_52_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17070_ clknet_leaf_27_wb_clk_i _02757_ _01053_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10514_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[31\] net790 net768 _06837_
+ _06842_ vssd1 vssd1 vccd1 vccd1 _06854_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_21_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14282_ net1336 vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_21_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11494_ net367 _07774_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[16\] net875
+ vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_150_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13185__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16021_ net1328 vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__inv_2
X_13233_ net2697 net352 net348 team_01_WB.instance_to_wrap.cpu.f0.i\[17\] vssd1 vssd1
+ vccd1 vccd1 _01917_ sky130_fd_sc_hd__a22o_1
XANTENNA__11697__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12292__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10445_ net1147 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[26\] net946
+ vssd1 vssd1 vccd1 vccd1 _06785_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_94_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13164_ net111 net849 net841 net1764 vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__a22o_1
X_10376_ net1144 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[16\] net975
+ vssd1 vssd1 vccd1 vccd1 _06716_ sky130_fd_sc_hd__and3_1
XFILLER_0_131_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12115_ net2131 net302 net456 vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__mux2_1
XANTENNA__16061__Q team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17972__1487 vssd1 vssd1 vccd1 vccd1 _17972__1487/HI net1487 sky130_fd_sc_hd__conb_1
X_17972_ net1487 vssd1 vssd1 vccd1 vccd1 la_data_out[14] sky130_fd_sc_hd__buf_2
X_13095_ net66 net65 net68 net67 vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__or4_2
XANTENNA__13488__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16923_ clknet_leaf_73_wb_clk_i _02610_ _00906_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_12046_ net2354 net227 net464 vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__mux2_1
X_16854_ clknet_leaf_29_wb_clk_i _02541_ _00837_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_140_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10171__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15805_ net1199 vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16785_ clknet_leaf_115_wb_clk_i _02472_ _00768_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13997_ net1684 net604 _04288_ net1185 vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12948_ net357 _03707_ _03708_ net870 net1974 vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__a32o_1
X_15736_ net1212 vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09864__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13660__A1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15667_ net1393 vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__inv_2
X_12879_ net1861 net872 net359 _03660_ vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__a22o_1
XANTENNA__12467__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17406_ clknet_leaf_82_wb_clk_i _03093_ _01389_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14618_ net1325 vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15598_ net1294 vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10495__B net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17337_ clknet_leaf_71_wb_clk_i _03024_ _01320_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14549_ net1410 vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10777__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08070_ _04537_ _04546_ vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload101 clknet_leaf_133_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload101/Y sky130_fd_sc_hd__clkinv_8
X_17268_ clknet_leaf_20_wb_clk_i _02955_ _01251_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload112 clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload112/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_114_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload123 clknet_leaf_108_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload123/Y sky130_fd_sc_hd__clkinv_4
Xclkload134 clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload134/Y sky130_fd_sc_hd__inv_4
XFILLER_0_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload145 clknet_leaf_86_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload145/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_114_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16219_ clknet_leaf_140_wb_clk_i net1614 _00207_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__dfrtp_1
X_17199_ clknet_leaf_33_wb_clk_i _02886_ _01182_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10529__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12923__B1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09508__C net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10934__C1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08412__C net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15807__A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08972_ net1007 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[8\] net896 vssd1
+ vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__and3_1
XFILLER_0_53_5 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09364__X _05704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09147__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold18 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[1\] vssd1 vssd1 vccd1 vccd1
+ net1553 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14140__A2 _04241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold29 team_01_WB.instance_to_wrap.cpu.f0.write_data\[4\] vssd1 vssd1 vccd1 vccd1
+ net1564 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08355__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout364_A _03580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09524_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[29\] net783 _05861_ _05862_
+ _05863_ vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_78_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09855__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09540__A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09455_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[29\] net694 _05792_
+ _05793_ _05794_ vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_78_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12377__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout531_A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1273_A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08406_ _04741_ _04744_ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13403__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09386_ _05713_ _05718_ _05725_ net703 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__o32a_4
XFILLER_0_4_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08337_ net1131 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[30\] net954
+ vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1061_X net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout417_X net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08268_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[13\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[5\]
+ net1050 vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout998_A _04491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08199_ net2448 net2359 net1052 vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__mux2_1
XANTENNA__12914__B1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10230_ net1143 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[9\] net977 vssd1
+ vssd1 vccd1 vccd1 _06570_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_35_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout786_X net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08594__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10161_ _06499_ _06500_ vssd1 vssd1 vccd1 vccd1 _06501_ sky130_fd_sc_hd__nor2_1
XANTENNA__12840__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1005 net1015 vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1016 net1031 vssd1 vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__clkbuf_4
Xfanout1027 net1028 vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__clkbuf_2
X_10092_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[7\] net804 net756 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06432_ sky130_fd_sc_hd__a22o_1
Xfanout1038 net1041 vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__buf_2
XANTENNA_fanout953_X net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17705__Q team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1049 net1059 vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__clkbuf_2
X_13920_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[12\] _04142_ _04207_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__a31o_1
X_13851_ net1180 net1067 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[12\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[12\] sky130_fd_sc_hd__and3b_1
XFILLER_0_88_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12802_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] net1062 net364 _03629_
+ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__a22o_1
XANTENNA__15452__A net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13782_ _04162_ _04165_ vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_48_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16570_ clknet_leaf_143_wb_clk_i _02257_ _00553_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11102__C1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10994_ _06399_ _07010_ vssd1 vssd1 vccd1 vccd1 _07334_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_48_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08992__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09310__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12733_ net1061 team_01_WB.instance_to_wrap.cpu.RU0.state\[0\] net638 vssd1 vssd1
+ vccd1 vccd1 _03583_ sky130_fd_sc_hd__o21ba_2
X_15521_ net1283 vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__inv_2
XANTENNA__12287__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11653__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15452_ net1245 vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_26_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ net2083 net202 net387 vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__mux2_1
X_14403_ net1360 vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11615_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] _07820_ vssd1 vssd1
+ vccd1 vccd1 _07830_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_137_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_74_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15383_ net1249 vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_96_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12595_ net2973 net208 net397 vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17122_ clknet_leaf_75_wb_clk_i _02809_ _01105_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_14334_ net1333 vssd1 vssd1 vccd1 vccd1 _00128_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11546_ net1713 net1173 net590 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] vssd1
+ vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13158__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17053_ clknet_leaf_69_wb_clk_i _02740_ _01036_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_14265_ net1224 vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11477_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[24\] net580 vssd1 vssd1 vccd1
+ vccd1 _07766_ sky130_fd_sc_hd__nand2_1
XANTENNA__11708__A1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16004_ net1348 vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__inv_2
X_13216_ _04505_ team_01_WB.instance_to_wrap.cpu.f0.state\[6\] _07649_ vssd1 vssd1
+ vccd1 vccd1 _03740_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_111_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09377__A2 _04808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10428_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[27\] net821 net749 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[27\]
+ _06767_ vssd1 vssd1 vccd1 vccd1 _06768_ sky130_fd_sc_hd__a221o_1
X_14196_ net1427 _04461_ _04462_ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_111_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13147_ net1693 net850 net842 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[29\] vssd1
+ vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__a22o_1
X_10359_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[17\] net776 net774 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _06699_ sky130_fd_sc_hd__a22o_1
XANTENNA__10392__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09625__A net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14122__A2 _04226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17955_ net1470 vssd1 vssd1 vccd1 vccd1 irq[0] sky130_fd_sc_hd__buf_2
XFILLER_0_57_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13078_ net3069 net2750 net852 vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__mux2_1
XANTENNA__13851__A_N net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12029_ net2540 net214 net465 vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__mux2_1
X_16906_ clknet_leaf_30_wb_clk_i _02593_ _00889_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_17886_ net107 vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10144__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10695__A1 _06902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16837_ clknet_leaf_47_wb_clk_i _02524_ _00820_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_109_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09063__C net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16768_ clknet_leaf_48_wb_clk_i _02455_ _00751_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13633__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15719_ net1389 vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__inv_2
XANTENNA__11644__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12197__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16699_ clknet_leaf_74_wb_clk_i _02386_ _00682_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_09240_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[21\] net677 net653 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[21\]
+ _05579_ vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09171_ net1010 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[16\] net934 vssd1
+ vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12925__S net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08122_ _04497_ team_01_WB.instance_to_wrap.cpu.f0.i\[3\] _04468_ team_01_WB.instance_to_wrap.cpu.f0.num\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_wire966_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08812__A1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08704__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13149__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08053_ _04512_ _04527_ vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08423__B net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09368__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09222__D1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_131_Right_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08040__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12660__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1021_A net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10383__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire921_X net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_119_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09535__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08955_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[6\] net668 _05278_ _05280_
+ _05286_ vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__a2111o_1
XANTENNA__14113__A2 _04265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout481_A _07949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout579_A _07752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08886_ net1107 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[2\] net915 vssd1
+ vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__and3_1
XANTENNA__10135__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08879__B2 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_16_Left_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10968__X _07308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12896__A _04837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout746_A net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15272__A net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09828__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08438__X _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09507_ net1150 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[29\] net974
+ vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout534_X net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09701__C net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09438_ _05764_ _05765_ _05776_ _05777_ vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__or4_1
XFILLER_0_94_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17971__1486 vssd1 vssd1 vccd1 vccd1 _17971__1486/HI net1486 sky130_fd_sc_hd__conb_1
XFILLER_0_149_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout701_X net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09369_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[26\] _04766_ net685
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[26\] _05708_ vssd1 vssd1 vccd1
+ vccd1 _05709_ sky130_fd_sc_hd__a221o_1
XFILLER_0_81_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12835__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11400_ _04469_ _07723_ _07721_ vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12380_ net2509 net280 net424 vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_25_Left_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11331_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[3\] net1176 _04552_ _07652_ vssd1
+ vssd1 vccd1 vccd1 _07664_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_158_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08333__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14054__C _04258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09359__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14050_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[43\] _04256_ _04262_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[51\]
+ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11262_ _06135_ _06163_ _07175_ net563 vssd1 vssd1 vccd1 vccd1 _07602_ sky130_fd_sc_hd__o31ai_1
X_13001_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[85\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[93\]
+ net859 vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__mux2_1
X_10213_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[8\] net797 net772 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _06553_ sky130_fd_sc_hd__a22o_1
XANTENNA__13560__B1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12570__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08031__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11193_ _07532_ net562 _07112_ vssd1 vssd1 vccd1 vccd1 _07533_ sky130_fd_sc_hd__and3b_1
XANTENNA__12423__X _03562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input42_A wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10144_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[11\] net821 net777 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06484_ sky130_fd_sc_hd__a22o_1
XANTENNA__14104__A2 _04236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17740_ clknet_leaf_92_wb_clk_i _03416_ _01680_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10075_ net1137 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[7\] net977 vssd1
+ vssd1 vccd1 vccd1 _06415_ sky130_fd_sc_hd__and3_1
X_14952_ net1375 vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_34_Left_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10126__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13903_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[4\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[6\] _04141_ vssd1 vssd1 vccd1 vccd1
+ _04204_ sky130_fd_sc_hd__and4_1
XANTENNA__10677__A1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17671_ clknet_leaf_0_wb_clk_i _03356_ _01612_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14883_ net1250 vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__inv_2
XANTENNA__11914__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16622_ clknet_leaf_28_wb_clk_i _02309_ _00605_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13834_ net1709 net830 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[27\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_134_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_139_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13765_ net1184 _04153_ vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__nand2_2
X_16553_ clknet_leaf_0_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[19\]
+ _00536_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13414__B _05224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10977_ net373 net341 net340 _06526_ net550 net539 vssd1 vssd1 vccd1 vccd1 _07317_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_104_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15504_ net1271 vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__inv_2
X_12716_ net2056 net306 net386 vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__mux2_1
X_13696_ _04502_ _04113_ _04117_ _04118_ vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__or4_2
X_16484_ clknet_leaf_152_wb_clk_i _02238_ _00467_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12647_ net2155 net297 net393 vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__mux2_1
X_15435_ net1423 vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_80_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15366_ net1383 vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_152_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12578_ net2950 net282 net399 vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_152_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08524__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17105_ clknet_leaf_112_wb_clk_i _02792_ _01088_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11529_ net1844 net1172 net588 net1080 vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__a22o_1
X_14317_ net1308 vssd1 vssd1 vccd1 vccd1 _00111_ sky130_fd_sc_hd__inv_2
X_15297_ net1278 vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__inv_2
Xhold307 team_01_WB.instance_to_wrap.a1.ADR_I\[23\] vssd1 vssd1 vccd1 vccd1 net1842
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10492__C net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold318 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1853 sky130_fd_sc_hd__dlygate4sd3_1
Xhold329 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1864 sky130_fd_sc_hd__dlygate4sd3_1
X_14248_ net1230 vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__inv_2
X_17036_ clknet_leaf_147_wb_clk_i _02723_ _01019_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09058__C net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12480__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14179_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[10\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[9\]
+ _04448_ vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__and3_1
Xfanout809 net810 vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08897__C net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09770__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08740_ net1017 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[4\] net902 vssd1
+ vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__and3_1
Xhold1007 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 net2542
+ sky130_fd_sc_hd__dlygate4sd3_1
X_17938_ net1453 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
Xhold1018 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[41\] vssd1 vssd1 vccd1 vccd1
+ net2553 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2564 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09522__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1380 net1384 vssd1 vssd1 vccd1 vccd1 net1380 sky130_fd_sc_hd__buf_2
Xfanout1391 net1398 vssd1 vssd1 vccd1 vccd1 net1391 sky130_fd_sc_hd__buf_2
X_08671_ net1006 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[7\] net923 vssd1
+ vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__and3_1
X_17869_ clknet_leaf_129_wb_clk_i _03544_ _01809_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_124_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08418__B net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09223_ _05554_ _05555_ _05556_ _05562_ vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__or4_1
XFILLER_0_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10840__A1 _06158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12655__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09154_ _04947_ _05492_ vssd1 vssd1 vccd1 vccd1 _05494_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08105_ team_01_WB.instance_to_wrap.cpu.f0.state\[2\] team_01_WB.instance_to_wrap.cpu.f0.state\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09085_ net1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[13\] net882
+ vssd1 vssd1 vccd1 vccd1 _05425_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09817__X _06157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08036_ net1744 net567 net345 team_01_WB.instance_to_wrap.cpu.f0.i\[19\] vssd1 vssd1
+ vccd1 vccd1 _03555_ sky130_fd_sc_hd__a22o_1
Xhold830 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold841 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold852 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2387 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout696_A _04766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold863 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[10\] vssd1 vssd1 vccd1 vccd1
+ net2398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold874 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold885 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2420 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1024_X net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1403_A net1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold896 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2431 sky130_fd_sc_hd__dlygate4sd3_1
X_09987_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[2\] net803 net758 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06327_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout484_X net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08938_ net1112 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[6\] net920 vssd1
+ vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__and3_1
XFILLER_0_99_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1530 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net3065 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10659__A1 _06188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1541 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net3076 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09513__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout651_X net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08869_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[3\] net657 _05191_ _05192_
+ _05201_ vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__a2111o_1
Xhold1552 _03486_ vssd1 vssd1 vccd1 vccd1 net3087 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_153_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1563 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net3098 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout749_X net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1574 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net3109 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08721__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10900_ net520 _06969_ _07236_ vssd1 vssd1 vccd1 vccd1 _07240_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_28_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1585 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[14\] vssd1 vssd1 vccd1 vccd1
+ net3120 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_28_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1596 team_01_WB.instance_to_wrap.cpu.K0.code\[6\] vssd1 vssd1 vccd1 vccd1 net3131
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11880_ net2786 net225 net483 vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__mux2_1
XANTENNA__11608__A0 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10831_ net562 _07089_ _07155_ _07170_ vssd1 vssd1 vccd1 vccd1 _07171_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_84_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout916_X net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13550_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] _05616_ _03925_ vssd1
+ vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10762_ _06945_ _07100_ net327 _06894_ vssd1 vssd1 vccd1 vccd1 _07102_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12501_ net2514 net270 net409 vssd1 vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__mux2_1
XANTENNA__10831__A1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13481_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] _05679_ _03941_ vssd1
+ vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12565__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10693_ _06889_ _06907_ net536 vssd1 vssd1 vccd1 vccd1 _07033_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15220_ net1378 vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__inv_2
X_12432_ net3112 net204 net415 vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15151_ net1300 vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_130_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12363_ net2064 net247 net425 vssd1 vssd1 vccd1 vccd1 _02633_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14102_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[93\] _04241_ _04262_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[53\]
+ _04388_ vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__a221o_1
X_11314_ team_01_WB.instance_to_wrap.cpu.f0.state\[3\] net1176 vssd1 vssd1 vccd1 vccd1
+ _07651_ sky130_fd_sc_hd__or2_1
X_15082_ net1283 vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__inv_2
X_12294_ net3049 net220 net433 vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14033_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[82\] _04245_ _04255_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[114\]
+ vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__a22o_1
XANTENNA__11909__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11245_ net523 _07248_ _07584_ vssd1 vssd1 vccd1 vccd1 _07585_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_121_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10898__A1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09752__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11176_ net525 _07158_ vssd1 vssd1 vccd1 vccd1 _07516_ sky130_fd_sc_hd__or2_1
XANTENNA__13409__B _05220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09606__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08510__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10127_ _05301_ _06466_ vssd1 vssd1 vccd1 vccd1 _06467_ sky130_fd_sc_hd__xor2_1
X_15984_ net1355 vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__inv_2
XANTENNA__09462__X _05802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17723_ clknet_leaf_156_wb_clk_i _00016_ _01664_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.state\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_145_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10058_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] net627 _06396_ _06397_
+ vssd1 vssd1 vccd1 vccd1 _06398_ sky130_fd_sc_hd__a22o_2
X_14935_ net1215 vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17654_ clknet_leaf_4_wb_clk_i net2011 _01595_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_14866_ net1290 vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__inv_2
XANTENNA__09114__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16605_ clknet_leaf_65_wb_clk_i _02292_ _00588_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13817_ net3075 net834 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[10\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_102_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17585_ clknet_leaf_124_wb_clk_i _03272_ _01544_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.code\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09268__A1 net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14797_ net1265 vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_69_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__15640__A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16536_ clknet_leaf_6_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[2\]
+ _00519_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_156_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13748_ team_01_WB.instance_to_wrap.cpu.c0.count\[3\] team_01_WB.instance_to_wrap.cpu.c0.count\[2\]
+ team_01_WB.instance_to_wrap.cpu.c0.count\[1\] vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_154_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12475__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16467_ clknet_leaf_12_wb_clk_i _02221_ _00450_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14256__A net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13679_ team_01_WB.instance_to_wrap.cpu.c0.count\[4\] team_01_WB.instance_to_wrap.cpu.c0.count\[5\]
+ _04101_ vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__and3_1
XANTENNA__08491__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15418_ net1370 vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__inv_2
X_16398_ clknet_leaf_93_wb_clk_i net1801 _00381_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15349_ net1275 vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__inv_2
XANTENNA__09440__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold104 net106 vssd1 vssd1 vccd1 vccd1 net1639 sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 _03527_ vssd1 vssd1 vccd1 vccd1 net1650 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09991__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold126 team_01_WB.instance_to_wrap.cpu.f0.write_data\[12\] vssd1 vssd1 vccd1 vccd1
+ net1661 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08541__X _04881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold137 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[122\] vssd1 vssd1 vccd1 vccd1
+ net1672 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11819__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13524__B1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold148 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[14\] vssd1 vssd1 vccd1 vccd1
+ net1683 sky130_fd_sc_hd__dlygate4sd3_1
X_17019_ clknet_leaf_71_wb_clk_i _02706_ _01002_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold159 _01995_ vssd1 vssd1 vccd1 vccd1 net1694 sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] net626 _06248_ _06249_
+ vssd1 vssd1 vccd1 vccd1 _06250_ sky130_fd_sc_hd__a22o_2
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout606 _03583_ vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__clkbuf_4
X_09841_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[13\] net819 net772 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06181_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09743__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout628 _03739_ vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkload14_A clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout639 _03572_ vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__clkbuf_2
X_17970__1485 vssd1 vssd1 vccd1 vccd1 _17970__1485/HI net1485 sky130_fd_sc_hd__conb_1
X_09772_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[15\] net822 net780 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_126_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08723_ net1097 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[5\] net919 vssd1
+ vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08703__B1 _05041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08654_ net1102 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[10\] net880
+ vssd1 vssd1 vccd1 vccd1 _04994_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_1_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08585_ net1104 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[15\] net890
+ vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout444_A _07959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15550__A net1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12802__A2 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12385__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10694__A _06906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout611_A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout232_X net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08435__Y _04775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1353_A net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09206_ net1005 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[17\] net878
+ vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09137_ net1022 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[14\] net907
+ vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1141_X net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09982__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09068_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[12\] net687 _05382_ _05400_
+ _05401_ vssd1 vssd1 vccd1 vccd1 _05408_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08451__X _04791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12318__A1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout699_X net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08019_ _04512_ _04514_ vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold660 team_01_WB.instance_to_wrap.cpu.RU0.state\[2\] vssd1 vssd1 vccd1 vccd1 net2195
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 _02064_ vssd1 vssd1 vccd1 vccd1 net2206 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12869__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11030_ _05455_ net373 vssd1 vssd1 vccd1 vccd1 _07370_ sky130_fd_sc_hd__and2_1
Xhold682 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2217 sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2228 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08330__C net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12981_ net2642 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[113\] net865 vssd1 vssd1
+ vccd1 vccd1 _02144_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_51_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1360 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2895 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1371 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[14\] vssd1 vssd1 vccd1 vccd1
+ net2906 sky130_fd_sc_hd__dlygate4sd3_1
X_14720_ net1187 vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__inv_2
Xhold1382 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 net2917
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11932_ net2639 net206 net477 vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1393 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[39\] vssd1 vssd1 vccd1 vccd1
+ net2928 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08339__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14651_ net1318 vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__inv_2
X_11863_ net2600 net215 net486 vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09161__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10814_ net343 _07091_ _07136_ _07153_ vssd1 vssd1 vccd1 vccd1 _07154_ sky130_fd_sc_hd__o31ai_4
X_13602_ net722 _07553_ net1076 vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__o21a_1
XFILLER_0_138_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17370_ clknet_leaf_76_wb_clk_i _03057_ _01353_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11794_ net3119 net220 net493 vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__mux2_1
X_14582_ net1401 vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16321_ clknet_leaf_119_wb_clk_i _02075_ _00304_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[44\]
+ sky130_fd_sc_hd__dfstp_1
X_10745_ _06906_ _07084_ net338 vssd1 vssd1 vccd1 vccd1 _07085_ sky130_fd_sc_hd__o21a_1
X_13533_ net196 net192 _07850_ net642 vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__o211a_1
XANTENNA__12295__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13464_ _03923_ _03924_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__and2_1
X_16252_ clknet_leaf_140_wb_clk_i net1730 _00240_ vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10280__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10676_ _07004_ _07015_ net529 vssd1 vssd1 vccd1 vccd1 _07016_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12415_ net2925 net278 net420 vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__mux2_1
XANTENNA__16064__Q team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15203_ net1234 vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__inv_2
XANTENNA__11212__B _07551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10568__A0 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13395_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] _04847_ vssd1 vssd1
+ vccd1 vccd1 _03856_ sky130_fd_sc_hd__xor2_1
X_16183_ clknet_leaf_7_wb_clk_i _01943_ _00171_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12346_ net2405 net251 net430 vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15134_ net1318 vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__inv_2
XANTENNA__09973__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_116_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_116_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15065_ net1238 vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__inv_2
X_12277_ net2279 net254 net436 vssd1 vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14016_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[65\] _04233_ _04245_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[81\]
+ _04306_ vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_75_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11228_ _06748_ _06749_ _05967_ vssd1 vssd1 vccd1 vccd1 _07568_ sky130_fd_sc_hd__a21o_1
XANTENNA__09725__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11159_ _06928_ _07497_ _07498_ _06920_ vssd1 vssd1 vccd1 vccd1 _07499_ sky130_fd_sc_hd__a22o_1
XANTENNA__09633__A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15967_ net1414 vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__inv_2
XANTENNA__10779__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17706_ clknet_leaf_134_wb_clk_i _03390_ _01647_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_14918_ net1404 vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15898_ net1352 vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_121_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17637_ clknet_leaf_157_wb_clk_i _03322_ _01578_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_148_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14849_ net1370 vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__inv_2
X_08370_ team_01_WB.instance_to_wrap.cpu.CU0.bit30 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\]
+ _04709_ vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__nand3_4
XFILLER_0_147_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17568_ clknet_leaf_87_wb_clk_i _03255_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16519_ clknet_leaf_0_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[17\]
+ _00502_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13993__B1 _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10718__S net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17499_ clknet_leaf_70_wb_clk_i _03186_ _01482_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12058__X _07955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10023__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11220__A1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09964__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11220__B2 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08431__B net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout403 net406 vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__buf_6
XANTENNA__09716__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout414 _03563_ vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__buf_4
Xfanout425 net426 vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__buf_6
Xfanout436 net438 vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13764__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09824_ _06159_ _06161_ vssd1 vssd1 vccd1 vccd1 _06164_ sky130_fd_sc_hd__xnor2_2
Xfanout447 _07958_ vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1101_A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout458 _07956_ vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__clkbuf_4
Xfanout469 net470 vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__clkbuf_8
Xclkbuf_4_14__f_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_14__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_09755_ _06073_ _06083_ _06084_ _06094_ vssd1 vssd1 vccd1 vccd1 _06095_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout659_A _04813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08706_ net1098 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[5\] net908 vssd1
+ vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__and3_1
X_09686_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[22\] net790 net730 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[22\]
+ _06003_ vssd1 vssd1 vccd1 vccd1 _06026_ sky130_fd_sc_hd__a221o_1
XANTENNA__08409__A_N _04738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08637_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[10\] net884 vssd1
+ vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_81_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout826_A _04579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout447_X net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08568_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[19\] net690 _04905_ _04906_
+ _04907_ vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_37_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12787__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13984__B1 _04258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout614_X net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10798__A0 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08499_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[3\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[2\]
+ _04622_ _04719_ vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__nand4_2
XFILLER_0_135_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10530_ _06865_ _06867_ _06869_ vssd1 vssd1 vccd1 vccd1 _06870_ sky130_fd_sc_hd__or3_1
XFILLER_0_92_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12539__A1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11032__B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10461_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[26\] net809 _06787_
+ _06791_ _06794_ vssd1 vssd1 vccd1 vccd1 _06801_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12843__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12200_ net2446 net201 net443 vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__mux2_1
XANTENNA__09277__X _05617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11211__A1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13180_ team_01_WB.instance_to_wrap.a1.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1
+ _03736_ sky130_fd_sc_hd__and2_1
X_10392_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[16\] net806 net742 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06732_ sky130_fd_sc_hd__a22o_1
X_12131_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[25\] net207 net453 vssd1
+ vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__mux2_1
X_12062_ net2537 net216 net461 vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__mux2_1
Xhold490 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[14\] vssd1 vssd1 vccd1 vccd1
+ net2025 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09156__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11013_ _07142_ _07143_ _07095_ vssd1 vssd1 vccd1 vccd1 _07353_ sky130_fd_sc_hd__a21boi_1
XPHY_EDGE_ROW_8_Left_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16870_ clknet_leaf_83_wb_clk_i _02557_ _00853_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout970 _04645_ vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_70_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15821_ net1192 vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__inv_2
Xfanout981 net983 vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_70_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout992 net993 vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__buf_2
XANTENNA__11194__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15752_ net1342 vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__inv_2
X_12964_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[0\] _05150_ net1039 vssd1
+ vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__mux2_1
XANTENNA__08143__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold1190 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[62\] vssd1 vssd1 vccd1 vccd1
+ net2725 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16059__Q team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14703_ net1198 vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__inv_2
X_11915_ net3148 net283 net482 vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__mux2_1
X_15683_ net1221 vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__inv_2
XANTENNA__08694__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12895_ net359 _03670_ _03671_ net872 net1589 vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__a32o_1
XANTENNA__11922__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17422_ clknet_leaf_37_wb_clk_i _03109_ _01405_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14634_ net1265 vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__inv_2
X_11846_ net3067 net286 net490 vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12778__A1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17353_ clknet_leaf_38_wb_clk_i _03040_ _01336_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11777_ net2235 net253 net495 vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14565_ net1410 vssd1 vssd1 vccd1 vccd1 _00359_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16304_ clknet_leaf_97_wb_clk_i _02058_ _00287_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10728_ net514 _07067_ vssd1 vssd1 vccd1 vccd1 _07068_ sky130_fd_sc_hd__nand2_1
X_13516_ net198 net194 _07837_ net644 vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__o211a_1
X_17284_ clknet_leaf_84_wb_clk_i _02971_ _01267_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_14496_ net1349 vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16235_ clknet_leaf_133_wb_clk_i net1694 _00223_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__dfrtp_1
X_13447_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] _05380_ vssd1 vssd1
+ vccd1 vccd1 _03908_ sky130_fd_sc_hd__xnor2_1
X_10659_ _06158_ _06188_ net546 vssd1 vssd1 vccd1 vccd1 _06999_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload13 clknet_leaf_156_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload13/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_77_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload24 clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload24/Y sky130_fd_sc_hd__bufinv_16
Xclkload35 clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload35/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_77_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload46 clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload46/Y sky130_fd_sc_hd__inv_8
XANTENNA__10005__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16166_ clknet_leaf_132_wb_clk_i _01929_ _00154_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13378_ _05834_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] vssd1 vssd1
+ vccd1 vccd1 _03839_ sky130_fd_sc_hd__and2b_1
Xclkload57 clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload57/Y sky130_fd_sc_hd__bufinv_16
Xclkload68 clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload68/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_149_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12950__A1 net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload79 clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload79/Y sky130_fd_sc_hd__inv_6
X_15117_ net1267 vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_114_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12329_ net2071 net211 net427 vssd1 vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16097_ clknet_leaf_115_wb_clk_i _01872_ _00085_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15048_ net1381 vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_3_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16999_ clknet_leaf_106_wb_clk_i _02686_ _00982_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_84_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09540_ net997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[28\] net949 vssd1
+ vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__and3_1
XANTENNA__13663__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_13_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09331__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09471_ net1002 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[30\] net918 vssd1
+ vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11832__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08422_ net1116 net1119 net1123 net1125 vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__and4b_1
XFILLER_0_59_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10956__B _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08353_ _04690_ _04691_ _04692_ vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__or3_1
XANTENNA__08426__B net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10244__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11441__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_74_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08284_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[3\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[2\]
+ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[1\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__and4b_1
XFILLER_0_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload7 clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload7/Y sky130_fd_sc_hd__inv_8
XFILLER_0_128_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12663__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout407_A _03564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1051_A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09398__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_25_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09538__A net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1316_A net1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14143__B1 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout200 _07858_ vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__buf_2
XANTENNA_fanout776_A _04667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1209 net1223 vssd1 vssd1 vccd1 vccd1 net1209 sky130_fd_sc_hd__buf_4
Xfanout211 net213 vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__buf_2
XANTENNA_fanout397_X net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout222 net224 vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__clkbuf_2
Xfanout233 net236 vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__buf_2
Xfanout244 _07862_ vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__clkbuf_2
Xfanout255 net256 vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1104_X net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout266 net268 vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__clkbuf_2
Xfanout277 net279 vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__clkbuf_2
X_09807_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[14\] net812 net780 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06147_ sky130_fd_sc_hd__a22o_1
Xfanout288 _07941_ vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__buf_2
Xfanout299 _07921_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__buf_1
X_07999_ team_01_WB.instance_to_wrap.cpu.f0.num\[3\] vssd1 vssd1 vccd1 vccd1 _04497_
+ sky130_fd_sc_hd__inv_2
XANTENNA_fanout943_A net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09704__C net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11308__A net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09738_ net1145 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[20\] net969
+ vssd1 vssd1 vccd1 vccd1 _06078_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09322__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11027__B _06158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout731_X net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12838__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09669_ net1144 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[22\] net951
+ vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__and3_1
XFILLER_0_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11742__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11700_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[11\] net717 vssd1 vssd1 vccd1
+ vccd1 _07897_ sky130_fd_sc_hd__or2_1
X_12680_ net2171 net298 net390 vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11631_ net2881 net245 net501 vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_64_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_148_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08336__B net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_145_Right_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10235__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14350_ net1333 vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__inv_2
XANTENNA__11432__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11562_ net3099 net1182 net35 vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13301_ net564 _03784_ net828 vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__a21o_1
X_10513_ _06849_ _06850_ _06851_ _06852_ vssd1 vssd1 vccd1 vccd1 _06853_ sky130_fd_sc_hd__or4_1
XFILLER_0_80_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14281_ net1336 vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12573__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10882__A _05566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11493_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[16\] net580 vssd1 vssd1 vccd1
+ vccd1 _07774_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_21_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13232_ net2900 net352 net348 team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1
+ vccd1 vccd1 _01918_ sky130_fd_sc_hd__a22o_1
X_16020_ net1328 vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__inv_2
XANTENNA__09928__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input72_A wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10444_ net1147 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[26\] net978
+ vssd1 vssd1 vccd1 vccd1 _06784_ sky130_fd_sc_hd__and3_1
XFILLER_0_150_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11196__A0 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10538__A3 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13163_ net1613 net851 net839 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[13\] vssd1
+ vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__a22o_1
X_10375_ _06712_ _06714_ vssd1 vssd1 vccd1 vccd1 _06715_ sky130_fd_sc_hd__nand2_1
XANTENNA__08600__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12114_ net2975 net281 net456 vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14134__B1 _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17971_ net1486 vssd1 vssd1 vccd1 vccd1 la_data_out[13] sky130_fd_sc_hd__buf_2
X_13094_ _03717_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[0\] net852 vssd1 vssd1
+ vccd1 vccd1 _02031_ sky130_fd_sc_hd__mux2_1
XANTENNA__11917__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16922_ clknet_leaf_76_wb_clk_i _02609_ _00905_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12045_ net2834 net286 net465 vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__mux2_1
XANTENNA__13417__B _05112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16853_ clknet_leaf_112_wb_clk_i _02540_ _00836_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15804_ net1199 vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__inv_2
X_16784_ clknet_leaf_144_wb_clk_i _02471_ _00767_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13996_ _04273_ _04275_ _04277_ _04287_ vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__or4_1
XFILLER_0_99_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09911__A _06250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15735_ net1244 vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__inv_2
X_12947_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[8\] net1039 vssd1 vssd1 vccd1
+ vccd1 _03708_ sky130_fd_sc_hd__or2_1
XANTENNA__11120__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13660__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11671__A1 _07232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15666_ net1267 vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__inv_2
X_12878_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[29\] _03659_ net1040 vssd1
+ vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__mux2_1
XANTENNA__08527__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17405_ clknet_leaf_65_wb_clk_i _03092_ _01388_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_14617_ net1308 vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11829_ net2190 net218 net489 vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__mux2_1
X_15597_ net1264 vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17336_ clknet_leaf_50_wb_clk_i _03023_ _01319_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14548_ net1407 vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10777__A3 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12483__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_131_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_131_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_17267_ clknet_leaf_24_wb_clk_i _02954_ _01250_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14264__A net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload102 clknet_leaf_134_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload102/X sky130_fd_sc_hd__clkbuf_4
X_14479_ net1399 vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__inv_2
Xclkload113 clknet_leaf_122_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload113/Y sky130_fd_sc_hd__inv_8
Xclkload124 clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload124/Y sky130_fd_sc_hd__bufinv_16
X_16218_ clknet_leaf_124_wb_clk_i net1765 _00206_ vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09919__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload135 clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload135/Y sky130_fd_sc_hd__inv_8
Xclkload146 clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload146/Y sky130_fd_sc_hd__inv_6
X_17198_ clknet_leaf_37_wb_clk_i _02885_ _01181_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16149_ clknet_leaf_128_wb_clk_i _01912_ _00137_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap967 _04650_ vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_87_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08971_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[8\] net693 _05308_ _05309_
+ _05310_ vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_121_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_109_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__17725__D net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11827__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold19 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[0\] vssd1 vssd1 vccd1 vccd1
+ net1554 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09093__A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09552__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09523_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[29\] net809 net746 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__a22o_1
XANTENNA__08658__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12658__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout357_A net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1099_A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09454_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[29\] net682 _04797_
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[29\] vssd1 vssd1 vccd1 vccd1
+ _05794_ sky130_fd_sc_hd__a22o_1
XANTENNA__11662__A1 _07135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08437__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08405_ _04732_ _04739_ _04740_ _04742_ vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__and4_1
XFILLER_0_143_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09385_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[26\] net647 _05720_
+ _05721_ _05724_ vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_108_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10217__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08336_ net1153 net955 vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08267_ net3120 net2352 net1042 vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__mux2_1
XANTENNA__12393__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_148_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_50_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08198_ net2407 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[75\] net1054 vssd1 vssd1
+ vccd1 vccd1 _03489_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout893_A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_89_Left_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12914__A1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08043__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1221_X net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14902__A net1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08594__A1 net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14116__B1 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10160_ net340 _06497_ _06498_ vssd1 vssd1 vccd1 vccd1 _06500_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout681_X net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout779_X net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1006 net1008 vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__buf_2
X_10091_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[7\] net817 net807 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06431_ sky130_fd_sc_hd__a22o_1
Xfanout1017 net1030 vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__buf_2
Xfanout1028 net1030 vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__buf_1
Xfanout1039 net1041 vssd1 vssd1 vccd1 vccd1 net1039 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout946_X net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13850_ net1179 net1066 net3182 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[11\]
+ sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_98_Left_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12801_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[9\] _07269_ net1035 vssd1 vssd1
+ vccd1 vccd1 _03629_ sky130_fd_sc_hd__mux2_1
XANTENNA__09731__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13781_ net1184 _04160_ _04163_ vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__and3_1
XANTENNA__10877__A net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10993_ net553 _07324_ _07332_ _07069_ vssd1 vssd1 vccd1 vccd1 _07333_ sky130_fd_sc_hd__o211ai_1
XANTENNA__12568__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15520_ net1272 vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__inv_2
XANTENNA__11653__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12732_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[31\] net1061 net362 _03581_
+ vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__a22o_1
XANTENNA__10456__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08347__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14068__B net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15451_ net1253 vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_26_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12663_ net2219 net204 net387 vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ net1356 vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__inv_2
XANTENNA__10208__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11614_ net719 _07056_ _07828_ vssd1 vssd1 vccd1 vccd1 _07829_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11405__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15382_ net1261 vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__inv_2
X_12594_ net2719 net247 net397 vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17121_ clknet_leaf_53_wb_clk_i _02808_ _01104_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14333_ net1338 vssd1 vssd1 vccd1 vccd1 _00127_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11545_ net1791 net1173 net590 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\] vssd1
+ vssd1 vccd1 vccd1 _03307_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_61_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17052_ clknet_leaf_50_wb_clk_i _02739_ _01035_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_14264_ net1226 vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__inv_2
X_11476_ net366 _07765_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[25\] net874
+ vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_151_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12905__A1 _03678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16003_ net1365 vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__inv_2
XANTENNA__08513__C net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08034__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13215_ net2 net836 net629 net1711 vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__o22a_1
X_10427_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[27\] net817 net755 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06767_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14195_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[16\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[15\]
+ _04458_ vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_111_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14812__A net1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10358_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[17\] net779 net749 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _06698_ sky130_fd_sc_hd__a22o_1
X_13146_ net1794 net850 net842 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[30\] vssd1
+ vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__a22o_1
XANTENNA__11647__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13077_ net2244 net2238 net866 vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__mux2_1
X_17954_ net1469 vssd1 vssd1 vccd1 vccd1 gpio_out[37] sky130_fd_sc_hd__buf_2
XFILLER_0_100_1006 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10289_ net1128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[19\] net956
+ vssd1 vssd1 vccd1 vccd1 _06629_ sky130_fd_sc_hd__and3_1
XANTENNA__13330__A1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16905_ clknet_leaf_39_wb_clk_i _02592_ _00888_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12028_ net2358 net219 net465 vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__mux2_1
X_17885_ clknet_leaf_135_wb_clk_i _03560_ _01825_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09344__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10123__Y _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16836_ clknet_leaf_82_wb_clk_i _02523_ _00819_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_109_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12478__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16767_ clknet_leaf_43_wb_clk_i _02454_ _00750_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10787__A _04919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14259__A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13979_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[32\] _04221_ _04246_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[40\]
+ vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__a22o_1
X_15718_ net1382 vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__inv_2
X_16698_ clknet_leaf_78_wb_clk_i _02385_ _00681_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15649_ net1278 vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09170_ _05499_ _05503_ _05505_ _05509_ vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__or4_1
XFILLER_0_56_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09065__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08121_ _04469_ team_01_WB.instance_to_wrap.cpu.f0.num\[26\] team_01_WB.instance_to_wrap.cpu.f0.num\[18\]
+ _04476_ vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__o22a_1
XFILLER_0_43_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17319_ clknet_leaf_107_wb_clk_i _03006_ _01302_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08812__A2 _05150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08052_ _04528_ _04529_ _04527_ vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_142_954 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10027__A net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09773__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08954_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[6\] net683 _05283_ _05285_
+ _05288_ vssd1 vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout1014_A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13321__A1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08885_ net1108 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[2\] net880 vssd1
+ vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout474_A _07952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12896__B net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13085__A0 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout641_A _03572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12388__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1383_A net1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout739_A net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09506_ net1150 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[29\] net976
+ vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__and3_1
XANTENNA__10438__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12832__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09437_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[28\] net681 net672 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[28\]
+ _05761_ vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_23_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout527_X net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout906_A _04785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1269_X net1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08454__X _04794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09368_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[26\] net681 net660 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08319_ net1139 net956 vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__and2_4
X_09299_ net1009 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[22\] net940 vssd1
+ vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__and3_1
XANTENNA_60 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11330_ _07663_ net1538 _07655_ vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout896_X net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11261_ _06163_ _07175_ _06135_ vssd1 vssd1 vccd1 vccd1 _07601_ sky130_fd_sc_hd__o21a_1
XANTENNA__14054__D _04259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12851__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12899__B1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10212_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[8\] net818 net808 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[8\]
+ _06551_ vssd1 vssd1 vccd1 vccd1 _06552_ sky130_fd_sc_hd__a221o_1
XANTENNA__13560__A1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13000_ net2878 net2841 net854 vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__mux2_1
X_11192_ _06598_ _06604_ _06742_ vssd1 vssd1 vccd1 vccd1 _07532_ sky130_fd_sc_hd__and3_1
XANTENNA__08630__A net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10143_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[11\] net811 net749 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06483_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13312__A1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09516__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14951_ net1396 vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__inv_2
X_10074_ net991 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[7\] net984 vssd1
+ vssd1 vccd1 vccd1 _06414_ sky130_fd_sc_hd__and3_1
XANTENNA_input35_A gpio_in[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09164__C net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13902_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[4\]
+ _04141_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[6\] vssd1 vssd1 vccd1 vccd1
+ _04203_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_89_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17670_ clknet_leaf_0_wb_clk_i _03355_ _01611_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14882_ net1320 vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__inv_2
XANTENNA__10103__C net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16621_ clknet_leaf_107_wb_clk_i _02308_ _00604_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13833_ net2115 net830 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[26\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__12298__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16552_ clknet_leaf_0_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[18\]
+ _00535_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11626__A1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10429__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13764_ team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[5\]
+ net604 vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__mux2_1
XANTENNA__10400__A net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10976_ _07015_ _07101_ _07312_ _07315_ vssd1 vssd1 vccd1 vccd1 _07316_ sky130_fd_sc_hd__a22o_1
X_17939__1454 vssd1 vssd1 vccd1 vccd1 _17939__1454/HI net1454 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_104_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15503_ net1388 vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_104_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12715_ net2138 net309 net384 vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__mux2_1
XANTENNA__08508__C net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16483_ clknet_leaf_140_wb_clk_i _02237_ _00466_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13695_ team_01_WB.instance_to_wrap.cpu.c0.count\[11\] team_01_WB.instance_to_wrap.cpu.c0.count\[8\]
+ team_01_WB.instance_to_wrap.cpu.c0.count\[15\] team_01_WB.instance_to_wrap.cpu.c0.count\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__or4bb_1
XANTENNA__11930__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15434_ net1284 vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__inv_2
X_12646_ net2271 net276 net391 vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_156_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08364__X _04704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08805__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15365_ net1287 vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__inv_2
X_12577_ net2386 net249 net402 vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_152_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_152_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17104_ clknet_leaf_21_wb_clk_i _02791_ _01087_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14316_ net1323 vssd1 vssd1 vccd1 vccd1 _00110_ sky130_fd_sc_hd__inv_2
X_11528_ net1664 net1172 net588 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\] vssd1
+ vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__a22o_1
X_15296_ net1272 vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__inv_2
Xhold308 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1843 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold319 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1854 sky130_fd_sc_hd__dlygate4sd3_1
X_17035_ clknet_leaf_5_wb_clk_i _02722_ _01018_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15638__A net1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12761__S net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14247_ net1218 vssd1 vssd1 vccd1 vccd1 _00041_ sky130_fd_sc_hd__inv_2
X_11459_ _04753_ _07630_ vssd1 vssd1 vccd1 vccd1 _07755_ sky130_fd_sc_hd__nor2_1
XANTENNA__08811__Y _05151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09636__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14178_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[9\] _04448_ net1996 vssd1
+ vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17626__Q team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13129_ net80 net846 net633 net1729 vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__a22o_1
XANTENNA__13303__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold1008 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2543 sky130_fd_sc_hd__dlygate4sd3_1
X_17937_ net1452 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
Xhold1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2554 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_128_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1370 net1373 vssd1 vssd1 vccd1 vccd1 net1370 sky130_fd_sc_hd__buf_4
X_08670_ net1086 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[7\] net929 vssd1
+ vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_128_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1381 net1383 vssd1 vssd1 vccd1 vccd1 net1381 sky130_fd_sc_hd__buf_4
X_17868_ clknet_leaf_127_wb_clk_i _03543_ _01808_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10668__A2 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1392 net1393 vssd1 vssd1 vccd1 vccd1 net1392 sky130_fd_sc_hd__buf_4
XFILLER_0_75_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16819_ clknet_leaf_24_wb_clk_i _02506_ _00802_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_17799_ clknet_leaf_100_wb_clk_i _03475_ _01739_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[69\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_124_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12001__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13180__X _03736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11840__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09222_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[17\] net690 _05544_ _05545_
+ net708 vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_17_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10840__A2 _06707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14031__A2 _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09153_ _04947_ _05492_ vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__and2_1
XANTENNA__12042__A1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08104_ team_01_WB.instance_to_wrap.cpu.f0.state\[2\] _04563_ _04574_ vssd1 vssd1
+ vccd1 vccd1 _04575_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10053__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09994__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09084_ net1012 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[13\] net905
+ vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13767__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08035_ net1826 net567 net345 team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1
+ vccd1 vccd1 _03556_ sky130_fd_sc_hd__a22o_1
Xhold820 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2355 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12671__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1131_A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold831 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2366 sky130_fd_sc_hd__dlygate4sd3_1
Xhold842 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2377 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13542__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1229_A net1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold853 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[40\] vssd1 vssd1 vccd1 vccd1
+ net2388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold864 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold875 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2410 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08450__A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11553__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout689_A _04773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold886 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2421 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold897 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[66\] vssd1 vssd1 vccd1 vccd1
+ net2432 sky130_fd_sc_hd__dlygate4sd3_1
X_09986_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[2\] net743 net771 vssd1
+ vssd1 vccd1 vccd1 _06326_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout1017_X net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08937_ net1028 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[6\] net942 vssd1
+ vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__and3_1
XANTENNA__11305__B1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout477_X net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1520 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net3055 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15283__A net1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1531 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net3066 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1542 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net3077 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08449__X _04789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08868_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[3\] net700 net679 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__a22o_1
Xhold1553 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net3088 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1564 team_01_WB.instance_to_wrap.cpu.K0.code\[5\] vssd1 vssd1 vccd1 vccd1 net3099
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1575 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net3110 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_28_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1586 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net3121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1597 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net3132 sky130_fd_sc_hd__dlygate4sd3_1
X_08799_ net1009 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[0\] net939 vssd1
+ vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout644_X net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10830_ _07169_ _07163_ _07162_ vssd1 vssd1 vccd1 vccd1 _07170_ sky130_fd_sc_hd__or3b_1
XANTENNA__11608__A1 _07019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12805__B1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08328__C net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12281__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10761_ net532 _06904_ vssd1 vssd1 vccd1 vccd1 _07101_ sky130_fd_sc_hd__nor2_1
XANTENNA__12846__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout811_X net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11750__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12820__A3 _03642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout909_X net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12500_ net2383 net244 net409 vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__mux2_1
XANTENNA__09029__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10692_ net533 _06896_ _07031_ net375 vssd1 vssd1 vccd1 vccd1 _07032_ sky130_fd_sc_hd__o211a_1
X_13480_ _03934_ _03936_ _03938_ _03940_ vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__o31a_1
XANTENNA__14022__A2 _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12431_ net2385 net274 net417 vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__mux2_1
XANTENNA__08344__B net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15150_ net1297 vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__inv_2
XANTENNA__09985__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12362_ net2596 net211 net423 vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14101_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[69\] _04247_ _04258_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[61\]
+ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11313_ _04504_ team_01_WB.instance_to_wrap.cpu.f0.state\[3\] net586 vssd1 vssd1
+ vccd1 vccd1 _00019_ sky130_fd_sc_hd__a21o_1
XANTENNA__12581__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15081_ net1293 vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__inv_2
X_12293_ net2570 net222 net431 vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08631__Y _04971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14032_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[42\] _04246_ _04263_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[122\]
+ _04312_ vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__a221o_1
X_11244_ _06906_ _06987_ _06991_ _05263_ _06903_ vssd1 vssd1 vccd1 vccd1 _07584_ sky130_fd_sc_hd__o221a_1
XFILLER_0_31_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11544__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11175_ net375 _06922_ _07068_ net528 vssd1 vssd1 vccd1 vccd1 _07515_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_56_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08960__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10126_ _05264_ _05265_ net377 vssd1 vssd1 vccd1 vccd1 _06466_ sky130_fd_sc_hd__o21ai_1
XANTENNA_input38_X net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1056 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15983_ net1413 vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__inv_2
XANTENNA__10418__A_N net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17722_ clknet_leaf_156_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_write_i
+ _01663_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.WRITE_I sky130_fd_sc_hd__dfrtp_2
X_14934_ net1261 vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__inv_2
X_10057_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[0\] net763 net622 vssd1
+ vssd1 vccd1 vccd1 _06397_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_106_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09191__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17653_ clknet_leaf_4_wb_clk_i _03338_ _01594_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14865_ net1423 vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__inv_2
XANTENNA_clkload0_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16604_ clknet_leaf_59_wb_clk_i _02291_ _00587_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13816_ net2077 net832 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[9\]
+ sky130_fd_sc_hd__and2_1
X_17584_ clknet_leaf_124_wb_clk_i _03271_ _01543_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.code\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10130__A _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14796_ net1258 vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16535_ clknet_leaf_6_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[1\]
+ _00518_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_13747_ _04504_ net3163 _07783_ team_01_WB.instance_to_wrap.cpu.DM0.state\[0\] vssd1
+ vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__a22o_1
X_10959_ _06958_ net327 _07295_ _07298_ vssd1 vssd1 vccd1 vccd1 _07299_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_154_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10283__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16466_ clknet_leaf_111_wb_clk_i _02220_ _00449_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13678_ team_01_WB.instance_to_wrap.cpu.c0.count\[3\] team_01_WB.instance_to_wrap.cpu.c0.count\[2\]
+ team_01_WB.instance_to_wrap.cpu.c0.count\[1\] team_01_WB.instance_to_wrap.cpu.c0.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__and4_1
XANTENNA__14013__A2 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_2__f_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15417_ net1239 vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__inv_2
X_12629_ net2741 net273 net392 vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16397_ clknet_leaf_122_wb_clk_i net1982 _00380_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_38_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15348_ net1400 vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10586__A1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15368__A net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold105 _02007_ vssd1 vssd1 vccd1 vccd1 net1640 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12491__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15279_ net1388 vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold116 net102 vssd1 vssd1 vccd1 vccd1 net1651 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[12\] vssd1 vssd1 vccd1 vccd1
+ net1662 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 _03528_ vssd1 vssd1 vccd1 vccd1 net1673 sky130_fd_sc_hd__dlygate4sd3_1
X_17018_ clknet_leaf_80_wb_clk_i _02705_ _01001_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09366__A net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13524__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold149 net158 vssd1 vssd1 vccd1 vccd1 net1684 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09840_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[13\] net806 net776 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[13\]
+ _06179_ vssd1 vssd1 vccd1 vccd1 _06180_ sky130_fd_sc_hd__a221o_1
Xfanout607 _03583_ vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__clkbuf_2
Xfanout629 _03739_ vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_13__f_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_13__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09771_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[15\] net778 net761 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[15\]
+ _06108_ vssd1 vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11835__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08722_ net1098 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[5\] net889 vssd1
+ vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08703__A1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08653_ net1102 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[10\] net919
+ vssd1 vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__and3_1
XANTENNA__09532__C net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09259__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08584_ net1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[15\] net920 vssd1
+ vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12263__A1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13864__A_N net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12666__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1081_A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout437_A net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13351__A team_01_WB.instance_to_wrap.cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1179_A net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14004__A2 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09205_ net1085 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[17\] net878
+ vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__and3_1
XFILLER_0_146_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13212__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10026__A0 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09136_ net1023 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[14\] net941 vssd1
+ vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__and3_1
XANTENNA__09967__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11223__C1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09431__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09067_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[12\] net693 _05390_ _05392_
+ _05398_ vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_8_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1134_X net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08018_ team_01_WB.instance_to_wrap.cpu.K0.code\[0\] _04513_ team_01_WB.instance_to_wrap.cpu.K0.code\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__or3b_2
XFILLER_0_103_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold650 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2185 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout973_A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09707__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold661 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2196 sky130_fd_sc_hd__dlygate4sd3_1
X_17938__1453 vssd1 vssd1 vccd1 vccd1 _17938__1453/HI net1453 sky130_fd_sc_hd__conb_1
XFILLER_0_124_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold672 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2207 sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2218 sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2229 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1301_X net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout761_X net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ _06305_ _06306_ _06307_ _06308_ vssd1 vssd1 vccd1 vccd1 _06309_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_86_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12980_ net2772 net2793 net863 vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_51_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1350 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2885 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1361 team_01_WB.instance_to_wrap.cpu.c0.count\[12\] vssd1 vssd1 vccd1 vccd1 net2896
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1372 team_01_WB.instance_to_wrap.cpu.f0.num\[9\] vssd1 vssd1 vccd1 vccd1 net2907
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11931_ net2084 net245 net477 vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__mux2_1
Xhold1383 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[62\] vssd1 vssd1 vccd1 vccd1
+ net2918 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1394 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2929 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11046__A net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14650_ net1240 vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__inv_2
X_11862_ net3029 net220 net485 vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13601_ net186 _04042_ _04043_ net725 vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__a211o_1
X_10813_ _07054_ _07151_ _07152_ _07148_ vssd1 vssd1 vccd1 vccd1 _07153_ sky130_fd_sc_hd__a211oi_4
X_14581_ net1414 vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12576__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11793_ net2147 net221 net491 vssd1 vssd1 vccd1 vccd1 _03181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16320_ clknet_leaf_95_wb_clk_i _02074_ _00303_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13532_ _03939_ _03940_ vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__xor2_1
X_10744_ _06986_ _06989_ net536 vssd1 vssd1 vccd1 vccd1 _07084_ sky130_fd_sc_hd__mux2_1
X_16251_ clknet_leaf_153_wb_clk_i net1576 _00239_ vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__dfrtp_1
X_13463_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] _05616_ vssd1 vssd1
+ vccd1 vccd1 _03924_ sky130_fd_sc_hd__xor2_1
XFILLER_0_129_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10675_ _07009_ _07014_ net517 vssd1 vssd1 vccd1 vccd1 _07015_ sky130_fd_sc_hd__mux2_2
X_15202_ net1316 vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__inv_2
X_12414_ net1864 net300 net420 vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16182_ clknet_leaf_7_wb_clk_i _01942_ _00170_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13394_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] _04885_ vssd1 vssd1
+ vccd1 vccd1 _03855_ sky130_fd_sc_hd__and2_1
XANTENNA__10568__A1 _06811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09422__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15133_ net1313 vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_58_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12345_ net2742 net227 net427 vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13506__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15064_ net1209 vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__inv_2
X_12276_ net3165 net259 net438 vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__mux2_1
XANTENNA__08090__A team_01_WB.instance_to_wrap.cpu.f0.i\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14015_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[65\] _04247_ _04265_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_75_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08521__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11227_ _06748_ _06749_ _05967_ vssd1 vssd1 vccd1 vccd1 _07567_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_75_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09914__A _06250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11158_ net530 _07049_ _07496_ vssd1 vssd1 vccd1 vccd1 _07498_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_156_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_156_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12880__B1_N net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10109_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[6\] net803 _04678_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06449_ sky130_fd_sc_hd__a22o_1
X_15966_ net1407 vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__inv_2
X_11089_ _07352_ _07422_ _07425_ _07341_ vssd1 vssd1 vccd1 vccd1 _07429_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09489__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14917_ net1286 vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__inv_2
X_17705_ clknet_leaf_134_wb_clk_i _03389_ _01646_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[26\]
+ sky130_fd_sc_hd__dfrtp_4
X_15897_ net1401 vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10498__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17636_ clknet_leaf_157_wb_clk_i _03321_ _01577_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_14848_ net1235 vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12486__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17567_ clknet_leaf_86_wb_clk_i _03254_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_14779_ net1250 vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16518_ clknet_leaf_1_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[16\]
+ _00501_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12796__A2 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17498_ clknet_leaf_77_wb_clk_i _03185_ _01481_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16449_ clknet_leaf_74_wb_clk_i _02203_ _00432_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10008__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10559__A1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09413__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Left_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout404 net406 vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__buf_6
Xfanout415 _03562_ vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__buf_8
Xfanout426 _07966_ vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__clkbuf_8
X_09823_ _06162_ vssd1 vssd1 vccd1 vccd1 _06163_ sky130_fd_sc_hd__inv_2
Xfanout437 net438 vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__buf_8
Xfanout448 _07958_ vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__buf_4
Xfanout459 _07955_ vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__buf_6
XANTENNA_fanout387_A _03569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09754_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[20\] net782 net759 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _06094_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08705_ net1017 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[5\] net881 vssd1
+ vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__and3_1
X_09685_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[22\] net814 net742 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[22\]
+ _06006_ vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_61_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1296_A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08636_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[10\] net893
+ vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_81_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10201__C net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13433__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout721_A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12396__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08567_ net999 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[19\] net891 vssd1
+ vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_54_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout819_A _04632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10247__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12787__A2 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10798__A1 _05898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08498_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[3\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[2\]
+ _04622_ _04719_ vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__and4_2
XFILLER_0_92_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09652__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09558__X _05898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10460_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[26\] net789 net731 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[26\]
+ _06799_ vssd1 vssd1 vccd1 vccd1 _06800_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_70_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08903__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11252__C_N net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09404__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09119_ net1023 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[14\] net916
+ vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10391_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[16\] net794 net733 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[16\]
+ _06717_ vssd1 vssd1 vccd1 vccd1 _06731_ sky130_fd_sc_hd__a221o_1
XANTENNA__08612__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_1__f_wb_clk_i_X clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12130_ net2934 net245 net453 vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout976_X net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08341__C net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12061_ net2622 net218 net461 vssd1 vssd1 vccd1 vccd1 _02924_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold480 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2015 sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 net2026
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11012_ _07341_ _07347_ _07349_ _07351_ vssd1 vssd1 vccd1 vccd1 _07352_ sky130_fd_sc_hd__nor4_1
XANTENNA__09734__A net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17724__Q team_01_WB.instance_to_wrap.cpu.RU0.state\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15820_ net1190 vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__inv_2
XANTENNA__13256__A team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout971 _04645_ vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout982 net983 vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout993 net994 vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10599__B _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_93_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15751_ net1341 vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_142_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09172__C net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11278__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12963_ net2101 net871 net358 _03716_ vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__a22o_1
XANTENNA__13672__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1180 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2715 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14702_ net1211 vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__inv_2
Xhold1191 _03468_ vssd1 vssd1 vccd1 vccd1 net2726 sky130_fd_sc_hd__dlygate4sd3_1
X_11914_ net2728 net249 net482 vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__mux2_1
X_15682_ net1321 vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12894_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[24\] net1040 vssd1 vssd1 vccd1
+ vccd1 _03671_ sky130_fd_sc_hd__or2_1
X_17421_ clknet_leaf_67_wb_clk_i _03108_ _01404_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_14633_ net1258 vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__inv_2
X_11845_ net1881 net253 net488 vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10238__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17352_ clknet_leaf_63_wb_clk_i _03039_ _01335_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_14564_ net1421 vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11776_ net3081 net259 net497 vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__mux2_1
XANTENNA__10789__A1 _04919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16303_ clknet_leaf_101_wb_clk_i net2308 _00286_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13515_ _03945_ _03947_ vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__xor2_1
XANTENNA__08516__C net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_109_Left_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10727_ _06968_ _07066_ net537 vssd1 vssd1 vccd1 vccd1 _07067_ sky130_fd_sc_hd__mux2_1
X_17283_ clknet_leaf_63_wb_clk_i _02970_ _01266_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_14495_ net1400 vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16234_ clknet_leaf_141_wb_clk_i net1617 _00222_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__dfrtp_1
X_13446_ _03905_ _03906_ vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__and2_1
X_10658_ _06216_ net340 net546 vssd1 vssd1 vccd1 vccd1 _06998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload14 clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload14/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload25 clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload25/Y sky130_fd_sc_hd__inv_6
X_16165_ clknet_leaf_134_wb_clk_i _01928_ _00153_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[28\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload36 clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload36/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_77_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload47 clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload47/Y sky130_fd_sc_hd__inv_8
X_13377_ net3090 net829 _03838_ team_01_WB.instance_to_wrap.cpu.f0.i\[0\] vssd1 vssd1
+ vccd1 vccd1 _01870_ sky130_fd_sc_hd__a22o_1
Xclkload58 clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload58/Y sky130_fd_sc_hd__clkinvlp_4
X_10589_ net375 _06928_ vssd1 vssd1 vccd1 vccd1 _06929_ sky130_fd_sc_hd__nand2_1
Xclkload69 clknet_leaf_52_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload69/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_149_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15116_ net1260 vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__inv_2
XANTENNA__12950__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12328_ net2809 net216 net429 vssd1 vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16096_ clknet_leaf_115_wb_clk_i _01871_ _00084_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_114_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15047_ net1389 vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12259_ net2020 net189 net435 vssd1 vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_118_Left_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16998_ clknet_leaf_83_wb_clk_i _02685_ _00981_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09082__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15949_ net1417 vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__inv_2
X_09470_ net1003 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[30\] net935 vssd1
+ vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08421_ net1002 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[23\] net940 vssd1
+ vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__and3_1
X_17619_ clknet_leaf_2_wb_clk_i _03304_ _01560_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10229__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11414__A team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_86_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_53_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_127_Left_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08352_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[30\] net791 net787 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__a22o_1
X_17937__1452 vssd1 vssd1 vccd1 vccd1 _17937__1452/HI net1452 sky130_fd_sc_hd__conb_1
XFILLER_0_11_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08283_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[1\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_138_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_27_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload8 clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload8/Y sky130_fd_sc_hd__inv_16
XANTENNA__09819__A _06158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08723__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10972__B net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13194__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13775__S net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_136_Left_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_1137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout201 net202 vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__buf_2
Xfanout212 net213 vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__buf_1
Xfanout223 net224 vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__buf_2
XANTENNA_fanout671_A _04797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout234 net236 vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__buf_2
Xfanout245 _07842_ vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__buf_2
XANTENNA_fanout769_A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout256 _07892_ vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__clkbuf_2
X_09806_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[14\] net783 net731 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06146_ sky130_fd_sc_hd__a22o_1
Xfanout267 net268 vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__buf_2
Xfanout278 net279 vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__buf_2
XANTENNA__10180__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout289 _07941_ vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__buf_1
X_07998_ team_01_WB.instance_to_wrap.cpu.f0.num\[6\] vssd1 vssd1 vccd1 vccd1 _04496_
+ sky130_fd_sc_hd__inv_2
X_09737_ net1132 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[20\] net984
+ vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout936_A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13654__B1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10468__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09668_ net994 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[22\] net956 vssd1
+ vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__and3_1
XANTENNA__08457__X _04797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08619_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[11\] net696 net656 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__a22o_1
XANTENNA__13406__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09599_ net996 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[24\] net952 vssd1
+ vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11324__A team_01_WB.instance_to_wrap.cpu.DM0.data_i\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11630_ _07839_ _07841_ net612 vssd1 vssd1 vccd1 vccd1 _07842_ sky130_fd_sc_hd__mux2_4
XFILLER_0_38_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11043__B _06250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11561_ net3131 net1182 net36 vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12854__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11611__X _07827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13300_ net1069 _07710_ vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_98_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10512_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[31\] net787 net730 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06852_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_98_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14280_ net1336 vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__inv_2
XANTENNA__08633__A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11492_ net367 _07773_ net2839 net874 vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_21_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09389__A1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13231_ net2680 net352 net348 team_01_WB.instance_to_wrap.cpu.f0.i\[19\] vssd1 vssd1
+ vccd1 vccd1 _01919_ sky130_fd_sc_hd__a22o_1
XANTENNA__13185__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10443_ net1147 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[26\] net949
+ vssd1 vssd1 vccd1 vccd1 _06783_ sky130_fd_sc_hd__and3b_1
XFILLER_0_122_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11196__A1 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08597__C1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input65_A wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13162_ net2142 net847 net839 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[14\] vssd1
+ vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__a22o_1
XANTENNA__09167__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10374_ _06713_ vssd1 vssd1 vccd1 vccd1 _06714_ sky130_fd_sc_hd__inv_2
XANTENNA__08920__X _05260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12113_ net3055 net251 net458 vssd1 vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17970_ net1485 vssd1 vssd1 vccd1 vccd1 la_data_out[12] sky130_fd_sc_hd__buf_2
X_13093_ _03716_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[1\] net852 vssd1 vssd1
+ vccd1 vccd1 _02032_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09464__A net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12044_ net1859 net254 net463 vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__mux2_1
X_16921_ clknet_leaf_104_wb_clk_i _02608_ _00904_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_144_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16852_ clknet_leaf_66_wb_clk_i _02539_ _00835_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10171__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout790 _04654_ vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__buf_6
X_15803_ net1217 vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__inv_2
X_16783_ clknet_leaf_28_wb_clk_i _02470_ _00766_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13995_ _04152_ _04283_ _04285_ _04286_ vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__or4_1
XANTENNA__11933__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15734_ net1269 vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__inv_2
XANTENNA__10459__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12946_ _05337_ _07757_ _03694_ vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_153_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09864__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15665_ net1398 vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__inv_2
X_12877_ _05802_ net577 net360 vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__o21ba_1
XANTENNA__09630__C net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17404_ clknet_leaf_58_wb_clk_i _03091_ _01387_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_14616_ net1310 vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__inv_2
X_11828_ net1761 net222 net487 vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__mux2_1
X_15596_ net1269 vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__inv_2
XANTENNA__14070__B1 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09616__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17335_ clknet_leaf_13_wb_clk_i _03022_ _01318_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_14547_ net1426 vssd1 vssd1 vccd1 vccd1 _00341_ sky130_fd_sc_hd__inv_2
XANTENNA__12764__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11759_ net1909 net189 net495 vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__mux2_1
XANTENNA__18017__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17266_ clknet_leaf_145_wb_clk_i _02953_ _01249_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09639__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14478_ net1350 vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_116_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload103 clknet_leaf_137_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload103/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_24_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16217_ clknet_leaf_124_wb_clk_i _01977_ _00205_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dfrtp_1
Xclkload114 clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload114/Y sky130_fd_sc_hd__clkinv_4
Xclkload125 clknet_leaf_73_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload125/Y sky130_fd_sc_hd__bufinv_16
X_13429_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\]
+ net595 vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17197_ clknet_leaf_67_wb_clk_i _02884_ _01180_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload136 clknet_leaf_95_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload136/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload147 clknet_leaf_89_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload147/Y sky130_fd_sc_hd__inv_6
XFILLER_0_23_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13581__C1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12923__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16148_ clknet_leaf_128_wb_clk_i _01911_ _00136_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10934__A1 _05338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08970_ net1007 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[8\] net914 vssd1
+ vssd1 vccd1 vccd1 _05310_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16079_ clknet_leaf_130_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[1\]
+ _00067_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[1\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_100_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_11_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17677__CLK clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08355__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12004__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput1 ACK_I vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08107__A2 net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11843__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09522_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[29\] net789 net780 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08718__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09855__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09453_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[29\] net689 net666 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__a22o_1
XANTENNA__09540__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout252_A _07904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10870__A0 _06098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08404_ _04743_ vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__inv_2
X_09384_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[26\] net669 _05722_ _05723_
+ vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__a211o_1
XFILLER_0_93_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14061__B1 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08335_ net992 net977 vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__and2_4
XFILLER_0_35_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12674__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1161_A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout517_A net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08266_ net3139 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[7\] net1044 vssd1 vssd1
+ vccd1 vccd1 _03421_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08197_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[84\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[76\]
+ net1044 vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1426_A net1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_144_Left_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12914__A2 _03684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09240__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15286__A net1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1081 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10090_ _06421_ _06427_ _06428_ _06429_ vssd1 vssd1 vccd1 vccd1 _06430_ sky130_fd_sc_hd__or4_1
Xfanout1007 net1008 vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__clkbuf_2
Xfanout1018 net1030 vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__clkbuf_2
Xfanout1029 net1030 vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout674_X net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11319__A team_01_WB.instance_to_wrap.cpu.DM0.data_i\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10223__A _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout841_X net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12849__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11753__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout939_X net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11606__X _07823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12800_ net1630 net639 net607 _03628_ vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_153_Left_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13780_ _04164_ vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10992_ net531 _07286_ _07331_ net558 vssd1 vssd1 vccd1 vccd1 _07332_ sky130_fd_sc_hd__a211o_1
XANTENNA__08503__C1 _04841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11102__B2 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[31\] _06961_ net1032 vssd1 vssd1
+ vccd1 vccd1 _03581_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11653__A2 _07621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08347__B net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15450_ net1371 vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12662_ net2512 net273 net389 vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ net1360 vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__inv_2
X_11613_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[29\] net715 net616 vssd1 vssd1
+ vccd1 vccd1 _07828_ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15381_ net1277 vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__inv_2
XANTENNA__12584__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12593_ net2686 net211 net395 vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_137_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14365__A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17120_ clknet_leaf_45_wb_clk_i _02807_ _01103_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14332_ net1338 vssd1 vssd1 vccd1 vccd1 _00126_ sky130_fd_sc_hd__inv_2
X_11544_ net1869 net1173 net590 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\] vssd1
+ vssd1 vccd1 vccd1 _03308_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_61_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17051_ clknet_leaf_70_wb_clk_i _02738_ _01034_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_14263_ net1204 vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__inv_2
XANTENNA__11501__B _07756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11475_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[25\] net579 vssd1 vssd1 vccd1
+ vccd1 _07765_ sky130_fd_sc_hd__nand2_1
X_16002_ net1353 vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13214_ net13 net838 net630 net2542 vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__a22o_1
X_10426_ _06763_ _06764_ _06765_ vssd1 vssd1 vccd1 vccd1 _06766_ sky130_fd_sc_hd__or3_1
X_14194_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[15\] _04458_ net2202 vssd1
+ vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11928__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13145_ net1702 net850 net842 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[31\] vssd1
+ vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__a22o_1
X_10357_ _06693_ _06694_ _06695_ _06696_ vssd1 vssd1 vccd1 vccd1 _06697_ sky130_fd_sc_hd__or4_1
XFILLER_0_21_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10392__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13076_ net2398 net2307 net864 vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__mux2_1
X_17953_ net1468 vssd1 vssd1 vccd1 vccd1 gpio_out[36] sky130_fd_sc_hd__buf_2
X_17936__1451 vssd1 vssd1 vccd1 vccd1 _17936__1451/HI net1451 sky130_fd_sc_hd__conb_1
XANTENNA__09729__B1_N net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10288_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[19\] net811 net794 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _06628_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16904_ clknet_leaf_26_wb_clk_i _02591_ _00887_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_12027_ net1776 net224 net463 vssd1 vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__mux2_1
XANTENNA__10133__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17884_ clknet_leaf_135_wb_clk_i _03559_ _01824_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10144__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09922__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16835_ clknet_leaf_26_wb_clk_i _02522_ _00818_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_109_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13444__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16766_ clknet_leaf_79_wb_clk_i _02453_ _00749_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13978_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[96\] _04244_ _04249_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10787__B net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15717_ net1262 vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__inv_2
X_12929_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[14\] net1040 vssd1 vssd1 vccd1
+ vccd1 _03696_ sky130_fd_sc_hd__or2_1
XANTENNA__11644__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16697_ clknet_leaf_100_wb_clk_i _02384_ _00680_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15648_ net1239 vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__inv_2
XANTENNA__14043__B1 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12494__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15579_ net1274 vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08120_ _04471_ team_01_WB.instance_to_wrap.cpu.f0.num\[24\] _04495_ net1069 vssd1
+ vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__o2bb2a_1
X_17318_ clknet_leaf_90_wb_clk_i _03005_ _01301_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08704__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13149__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08051_ team_01_WB.instance_to_wrap.cpu.K0.code\[7\] team_01_WB.instance_to_wrap.cpu.K0.code\[6\]
+ team_01_WB.instance_to_wrap.cpu.K0.code\[5\] team_01_WB.instance_to_wrap.cpu.K0.code\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__or4b_2
X_17249_ clknet_leaf_57_wb_clk_i _02936_ _01232_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10308__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09656__X _05996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10907__A1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11838__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08576__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10742__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09816__B net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10383__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08953_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[6\] net679 _05267_ _05274_
+ _05275_ vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09535__C net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11139__A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08884_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\] net729 _05111_ net1121 vssd1
+ vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__a22oi_4
XANTENNA__10135__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1007_A net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12669__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout467_A net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09828__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09505_ net1148 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[29\] net981
+ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout634_A _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12832__B2 _03650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09436_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[28\] net659 _05775_
+ net706 vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__a211o_1
XFILLER_0_19_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14034__B1 _04254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout801_A _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09367_ net603 _05705_ _05706_ vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_43_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout422_X net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11602__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08318_ net1158 net1161 net1164 net1166 vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__and4_1
XFILLER_0_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09298_ net1005 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[22\] net925 vssd1
+ vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__and3_1
XANTENNA_50 _03654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_61 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08249_ net3026 net2816 net1046 vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1429_X net1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11260_ net343 _07567_ _07590_ _07599_ vssd1 vssd1 vccd1 vccd1 _07600_ sky130_fd_sc_hd__o31a_2
XTAP_TAPCELL_ROW_91_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12899__A1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08470__X _04810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout791_X net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout889_X net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10211_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[8\] net801 net744 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _06551_ sky130_fd_sc_hd__a22o_1
XANTENNA__13560__A2 _07171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11191_ _07191_ _07521_ _07530_ vssd1 vssd1 vccd1 vccd1 _07531_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10142_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[11\] net787 net768 vssd1
+ vssd1 vccd1 vccd1 _06482_ sky130_fd_sc_hd__a21o_1
X_10073_ net1138 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[7\] net963 vssd1
+ vssd1 vccd1 vccd1 _06413_ sky130_fd_sc_hd__and3_1
X_14950_ net1404 vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__inv_2
X_13901_ net571 _04202_ vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__and2_1
XANTENNA__09742__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input28_A DAT_I[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14881_ net1278 vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__inv_2
XANTENNA__12579__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17732__Q team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13832_ net1643 net831 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[25\]
+ sky130_fd_sc_hd__and2_1
X_16620_ clknet_leaf_19_wb_clk_i _02307_ _00603_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16551_ clknet_leaf_0_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[17\]
+ _00534_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09180__C net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13763_ net604 vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_139_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10975_ _05301_ net372 net333 _07314_ vssd1 vssd1 vccd1 vccd1 _07315_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_104_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15502_ net1297 vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__inv_2
X_12714_ net1990 net293 net386 vssd1 vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16482_ clknet_leaf_153_wb_clk_i _02236_ _00465_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14025__B1 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13694_ team_01_WB.instance_to_wrap.cpu.c0.count\[6\] _04116_ team_01_WB.instance_to_wrap.cpu.c0.count\[5\]
+ _04101_ vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__or4b_1
XFILLER_0_73_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15433_ net1296 vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__inv_2
X_12645_ net2722 net300 net391 vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_156_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10047__D1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15364_ net1219 vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_80_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09452__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12576_ net2735 net225 net400 vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_152_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17103_ clknet_leaf_34_wb_clk_i _02790_ _01086_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_14315_ net1323 vssd1 vssd1 vccd1 vccd1 _00109_ sky130_fd_sc_hd__inv_2
XANTENNA__08524__C net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11527_ net1590 net1171 net588 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] vssd1
+ vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__a22o_1
X_15295_ net1314 vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__inv_2
XANTENNA__14823__A net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10128__A net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17034_ clknet_leaf_31_wb_clk_i _02721_ _01017_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold309 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[24\] vssd1 vssd1 vccd1 vccd1
+ net1844 sky130_fd_sc_hd__dlygate4sd3_1
X_14246_ net1218 vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__inv_2
X_11458_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[31\] net579 vssd1 vssd1 vccd1
+ vccd1 _07754_ sky130_fd_sc_hd__nand2_1
XANTENNA__08821__A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10409_ _06107_ _06747_ _05999_ _06102_ _06103_ vssd1 vssd1 vccd1 vccd1 _06749_ sky130_fd_sc_hd__o2111a_1
X_14177_ net2921 _04448_ _04450_ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__o21a_1
XFILLER_0_22_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_4_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11389_ team_01_WB.instance_to_wrap.cpu.f0.i\[30\] _07696_ _07716_ vssd1 vssd1 vccd1
+ vccd1 _07718_ sky130_fd_sc_hd__and3_1
X_13128_ net1658 net843 net631 team_01_WB.instance_to_wrap.a1.ADR_I\[15\] vssd1 vssd1
+ vccd1 vccd1 _02013_ sky130_fd_sc_hd__a22o_1
Xclkbuf_4_12__f_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_12__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__15654__A net1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17936_ net1451 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
X_13059_ net2958 net2856 net861 vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__mux2_1
Xhold1009 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2544 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1360 net1362 vssd1 vssd1 vccd1 vccd1 net1360 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_128_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1371 net1373 vssd1 vssd1 vccd1 vccd1 net1371 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_128_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1382 net1383 vssd1 vssd1 vccd1 vccd1 net1382 sky130_fd_sc_hd__buf_2
X_17867_ clknet_leaf_125_wb_clk_i _03542_ _01807_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1393 net1394 vssd1 vssd1 vccd1 vccd1 net1393 sky130_fd_sc_hd__buf_4
XANTENNA__17642__Q team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08730__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16818_ clknet_leaf_110_wb_clk_i _02505_ _00801_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_17798_ clknet_leaf_99_wb_clk_i _03474_ _01738_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[68\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_16_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09090__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16749_ clknet_leaf_108_wb_clk_i _02436_ _00732_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_52 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14016__B1 _04245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09221_ _05557_ _05558_ _05559_ _05560_ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_17_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10840__A3 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09152_ _05416_ _05454_ _05491_ vssd1 vssd1 vccd1 vccd1 _05492_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08103_ _04568_ _04571_ _04572_ _04573_ vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__or4_4
XANTENNA__08434__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08797__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09083_ net1094 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[13\] net934
+ vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__and3_1
XANTENNA__12952__S net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12805__X _03632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout215_A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08034_ net1737 net568 net347 team_01_WB.instance_to_wrap.cpu.f0.i\[21\] vssd1 vssd1
+ vccd1 vccd1 _03557_ sky130_fd_sc_hd__a22o_1
XANTENNA__09386__X _05726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput70 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_31_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold810 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2345 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold821 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold832 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2367 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold843 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2378 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08549__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold854 _02079_ vssd1 vssd1 vccd1 vccd1 net2389 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10356__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold865 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[41\] vssd1 vssd1 vccd1 vccd1
+ net2400 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08450__B net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold876 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2411 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold887 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2422 sky130_fd_sc_hd__dlygate4sd3_1
Xhold898 _03472_ vssd1 vssd1 vccd1 vccd1 net2433 sky130_fd_sc_hd__dlygate4sd3_1
X_09985_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[2\] net810 net732 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06325_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08936_ net1027 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[6\] net899 vssd1
+ vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__and3_1
XANTENNA__10108__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11305__A1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1510 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net3045 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10204__C net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09562__A _05898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1521 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net3056 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1532 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net3067 sky130_fd_sc_hd__dlygate4sd3_1
X_08867_ net1017 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[3\] net931 vssd1
+ vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__and3_1
XANTENNA__12399__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout751_A net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout372_X net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1543 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3078 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1554 team_01_WB.instance_to_wrap.a1.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 net3089
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1565 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net3100 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout849_A net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08721__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1576 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net3111 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_28_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10501__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08798_ net1093 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[0\] net939 vssd1
+ vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_28_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1587 team_01_WB.instance_to_wrap.cpu.K0.code\[1\] vssd1 vssd1 vccd1 vccd1 net3122
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1598 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[6\] vssd1 vssd1 vccd1 vccd1 net3133
+ sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_8_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12805__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout637_X net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10816__A0 _05996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10760_ net522 _06904_ vssd1 vssd1 vccd1 vccd1 _07100_ sky130_fd_sc_hd__nor2_2
XANTENNA__14007__B1 _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09682__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08906__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09419_ _05758_ vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout804_X net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10691_ _05190_ _06908_ vssd1 vssd1 vccd1 vccd1 _07031_ sky130_fd_sc_hd__nand2_1
X_12430_ net3088 net208 net417 vssd1 vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13230__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11241__A0 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08788__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12361_ net2441 net215 net423 vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12862__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_130_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14100_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[13\] _04226_ _04259_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[21\]
+ _04386_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__a221o_1
X_11312_ net829 _07649_ vssd1 vssd1 vccd1 vccd1 _07650_ sky130_fd_sc_hd__or2_4
X_15080_ net1377 vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__inv_2
XANTENNA__09737__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12292_ net2302 net188 net431 vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__mux2_1
XANTENNA__08641__A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17727__Q team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14031_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[66\] _04247_ _04262_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[50\]
+ _04310_ vssd1 vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__a221o_1
X_11243_ _06966_ _07527_ _06964_ vssd1 vssd1 vccd1 vccd1 _07583_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13259__A team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12741__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11174_ net370 _07511_ _07513_ net341 _05417_ vssd1 vssd1 vccd1 vccd1 _07514_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_56_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08960__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10125_ net506 _06464_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] net626
+ vssd1 vssd1 vccd1 vccd1 _06465_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_98_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15982_ net1405 vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17721_ clknet_leaf_156_wb_clk_i _00015_ _01662_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09472__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10056_ _06384_ _06385_ _06390_ _06395_ vssd1 vssd1 vccd1 vccd1 _06396_ sky130_fd_sc_hd__or4_4
X_14933_ net1287 vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17652_ clknet_leaf_15_wb_clk_i _03337_ _01593_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12102__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10411__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14864_ net1274 vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__inv_2
X_16603_ clknet_leaf_70_wb_clk_i _02290_ _00586_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08519__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13815_ net3185 net834 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[8\]
+ sky130_fd_sc_hd__and2_1
X_14795_ net1395 vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__inv_2
X_17583_ clknet_leaf_94_wb_clk_i _03270_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.lcd_rs
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11941__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09268__A3 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10807__B1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13746_ team_01_WB.instance_to_wrap.cpu.RU0.state\[0\] _03579_ _04137_ team_01_WB.instance_to_wrap.cpu.RU0.next_dhit
+ net831 vssd1 vssd1 vccd1 vccd1 _00014_ sky130_fd_sc_hd__a311o_1
X_16534_ clknet_leaf_6_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[0\]
+ _00517_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_85_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10958_ _05042_ _06924_ _07297_ net368 vssd1 vssd1 vccd1 vccd1 _07298_ sky130_fd_sc_hd__o211a_1
XANTENNA__08816__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13441__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13677_ team_01_WB.instance_to_wrap.cpu.c0.count\[1\] team_01_WB.instance_to_wrap.cpu.c0.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16465_ clknet_leaf_20_wb_clk_i _02219_ _00448_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10889_ _07017_ _07217_ _07218_ _07100_ _07226_ vssd1 vssd1 vccd1 vccd1 _07229_ sky130_fd_sc_hd__a221o_1
XFILLER_0_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12628_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[25\] net207 net392 vssd1
+ vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__mux2_1
X_15416_ net1213 vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16396_ clknet_leaf_96_wb_clk_i net2851 _00379_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09425__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15347_ net1421 vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__inv_2
X_12559_ net2689 net216 net401 vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10586__A2 _06882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15278_ net1298 vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold106 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[20\] vssd1 vssd1 vccd1 vccd1 net1641
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold117 _02003_ vssd1 vssd1 vccd1 vccd1 net1652 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08551__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold128 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[22\] vssd1 vssd1 vccd1 vccd1 net1663
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 team_01_WB.instance_to_wrap.cpu.f0.write_data\[16\] vssd1 vssd1 vccd1 vccd1
+ net1674 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13524__A2 _07588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16541__Q team_01_WB.instance_to_wrap.cpu.DM0.data_i\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14229_ net3071 vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__clkbuf_1
X_17017_ clknet_leaf_102_wb_clk_i _02704_ _01000_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_78_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09366__B _05704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12732__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11535__B2 net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout608 _03583_ vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09085__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08951__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09770_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[15\] net816 net809 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06110_ sky130_fd_sc_hd__a22o_1
X_08721_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[5\] net698 net669 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__a22o_1
X_17919_ net1526 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
XANTENNA__11299__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1190 net1192 vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__buf_4
XANTENNA__08703__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12012__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08652_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[10\] net924
+ vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__and3_1
XANTENNA__10321__A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10510__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08429__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08583_ net1104 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[15\] net903
+ vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11851__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12799__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_44_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_48_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1074_A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09204_ net1085 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[17\] net934
+ vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10026__A1 _06365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13778__S net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09135_ net1110 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[14\] net943
+ vssd1 vssd1 vccd1 vccd1 _05475_ sky130_fd_sc_hd__and3_1
XANTENNA__12682__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1241_A net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1339_A net1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09066_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[12\] net670 _05389_ _05393_
+ _05397_ vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout799_A _04649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08017_ team_01_WB.instance_to_wrap.cpu.K0.code\[3\] team_01_WB.instance_to_wrap.cpu.K0.code\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold640 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2175 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold651 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2186 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1127_X net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11526__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold662 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[25\] vssd1 vssd1 vccd1 vccd1 net2197
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold673 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2208 sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2219 sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2230 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout587_X net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11168__A_N _07323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09968_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[3\] net761 net750 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06308_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_34_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08919_ net603 _05224_ vssd1 vssd1 vccd1 vccd1 _05259_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_86_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_83_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout754_X net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09899_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[5\] net812 _06227_ _06232_
+ _06233_ vssd1 vssd1 vccd1 vccd1 _06239_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_86_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1340 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[10\] vssd1 vssd1 vccd1 vccd1
+ net2875 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11930_ net2207 net212 net475 vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__mux2_1
Xhold1351 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2886 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1362 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[48\] vssd1 vssd1 vccd1 vccd1
+ net2897 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1373 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2908 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1384 _02101_ vssd1 vssd1 vccd1 vccd1 net2919 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1395 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2930 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08339__C net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11861_ net1882 net223 net483 vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__mux2_1
XANTENNA__12857__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13600_ net197 net193 _07891_ net643 vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__o211a_1
XANTENNA__11761__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10812_ net558 _07141_ _07017_ vssd1 vssd1 vccd1 vccd1 _07152_ sky130_fd_sc_hd__o21a_1
X_14580_ net1421 vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13451__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11792_ net3103 net188 net491 vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__mux2_1
XANTENNA__08636__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13451__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13531_ _03984_ _03985_ net1074 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\]
+ vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_149_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10743_ _06990_ _06994_ net536 vssd1 vssd1 vccd1 vccd1 _07083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16250_ clknet_leaf_152_wb_clk_i net1608 _00238_ vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__dfrtp_1
X_13462_ _03855_ _03921_ _03853_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__o21a_1
XFILLER_0_36_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10674_ _07011_ _07013_ net541 vssd1 vssd1 vccd1 vccd1 _07014_ sky130_fd_sc_hd__mux2_1
XANTENNA__09407__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15201_ net1278 vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__inv_2
X_12413_ net2192 net280 net420 vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__mux2_1
X_16181_ clknet_leaf_7_wb_clk_i _01941_ _00169_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13393_ _03853_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__inv_2
XANTENNA__12592__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15132_ net1243 vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__inv_2
X_12344_ net2284 net286 net430 vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08802__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13506__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15063_ net1220 vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__inv_2
X_12275_ net2549 net230 net437 vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__mux2_1
XANTENNA__11517__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14014_ _04301_ _04302_ _04303_ _04304_ vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__or4_1
XFILLER_0_121_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09186__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11226_ net563 _07556_ _07557_ _07565_ vssd1 vssd1 vccd1 vccd1 _07566_ sky130_fd_sc_hd__a31o_2
XTAP_TAPCELL_ROW_75_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11936__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11157_ net524 _07025_ _07496_ vssd1 vssd1 vccd1 vccd1 _07497_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10108_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[6\] net762 _06446_ _06447_
+ vssd1 vssd1 vccd1 vccd1 _06448_ sky130_fd_sc_hd__a211o_1
X_15965_ net1418 vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__inv_2
X_11088_ _07340_ _07427_ vssd1 vssd1 vccd1 vccd1 _07428_ sky130_fd_sc_hd__nand2_1
XANTENNA__09633__C net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17704_ clknet_leaf_133_wb_clk_i _03388_ _01645_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[25\]
+ sky130_fd_sc_hd__dfrtp_4
X_10039_ net1142 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[0\] net973 vssd1
+ vssd1 vccd1 vccd1 _06379_ sky130_fd_sc_hd__and3_1
X_14916_ net1230 vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09894__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15896_ net1351 vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17635_ clknet_leaf_157_wb_clk_i _03320_ _01576_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_121_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12767__S net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_125_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_125_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_14847_ net1312 vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_121_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11671__S net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17566_ clknet_leaf_86_wb_clk_i _03253_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_14778_ net1312 vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__inv_2
XANTENNA__09110__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16517_ clknet_leaf_1_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[15\]
+ _00500_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11453__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16536__Q team_01_WB.instance_to_wrap.cpu.DM0.data_i\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13729_ team_01_WB.instance_to_wrap.cpu.DM0.state\[1\] team_01_WB.instance_to_wrap.cpu.DM0.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__or2_1
XANTENNA__13993__A2 _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17497_ clknet_leaf_71_wb_clk_i _03184_ _01480_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_128_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_156_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16448_ clknet_leaf_25_wb_clk_i _02202_ _00431_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_144_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15379__A net1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11205__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16379_ clknet_leaf_119_wb_clk_i net2842 _00362_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08712__C net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12007__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10316__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09031__D1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout405 net406 vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__buf_4
Xfanout416 _03562_ vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11846__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09822_ _06159_ _06161_ vssd1 vssd1 vccd1 vccd1 _06162_ sky130_fd_sc_hd__or2_1
Xfanout427 _07965_ vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__buf_6
XANTENNA__12720__A3 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout438 _07963_ vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__buf_8
Xfanout449 _07958_ vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__clkbuf_8
X_09753_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[20\] net731 _06090_ _06091_
+ _06092_ vssd1 vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout282_A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08704_ net1097 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[5\] net916 vssd1
+ vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__and3_1
XANTENNA__13130__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09334__C1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09684_ _06020_ _06021_ _06022_ _06023_ vssd1 vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__or4_1
XFILLER_0_154_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08635_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[10\] net936 vssd1
+ vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__and3_1
XANTENNA__12677__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1289_A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08566_ net999 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[19\] net887 vssd1
+ vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__and3_1
XANTENNA__13433__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13984__A2 _04230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08497_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[23\] net701 _04834_ _04836_
+ vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__o22a_4
XANTENNA_fanout714_A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout335_X net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10798__A2 _06779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1077_X net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13197__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout502_X net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09118_ net1023 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[14\] net880
+ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10390_ _06718_ _06721_ _06726_ _06729_ vssd1 vssd1 vccd1 vccd1 _06730_ sky130_fd_sc_hd__or4_1
X_09049_ net1029 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[12\] net937 vssd1
+ vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__and3_1
XANTENNA__10226__A _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12060_ net2536 net221 net459 vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__mux2_1
Xhold470 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2005 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold481 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2016 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout871_X net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08376__B1 _04710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout969_X net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11756__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11011_ _05681_ net511 vssd1 vssd1 vccd1 vccd1 _07351_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_53_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold492 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2027 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08915__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout950 _04665_ vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout972 net974 vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout994 net995 vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13121__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09876__A0 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15750_ net1342 vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__inv_2
X_12962_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[1\] _05187_ net1039 vssd1
+ vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_142_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08918__X _05258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1170 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2705 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input10_A DAT_I[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1181 team_01_WB.instance_to_wrap.cpu.f0.num\[1\] vssd1 vssd1 vccd1 vccd1 net2716
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14701_ net1211 vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__inv_2
X_11913_ net2916 net226 net479 vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__mux2_1
Xhold1192 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2727 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12587__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10896__A net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12893_ net361 _03669_ net1036 vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__o21ai_1
X_15681_ net1280 vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__inv_2
X_17420_ clknet_leaf_148_wb_clk_i _03107_ _01403_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_14632_ net1395 vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__inv_2
X_11844_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[14\] net260 net489 vssd1
+ vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__mux2_1
XANTENNA__09628__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14563_ net1427 vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17351_ clknet_leaf_105_wb_clk_i _03038_ _01334_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11775_ net2704 net231 net496 vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16302_ clknet_leaf_93_wb_clk_i _02056_ _00285_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10726_ _05867_ _05898_ net548 vssd1 vssd1 vccd1 vccd1 _07066_ sky130_fd_sc_hd__mux2_1
X_13514_ net988 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] _03970_ _03971_
+ vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__a22o_1
X_17282_ clknet_leaf_56_wb_clk_i _02969_ _01265_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_14494_ net1354 vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_836 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13188__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16233_ clknet_leaf_135_wb_clk_i net1679 _00221_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__dfrtp_1
X_13445_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] _05419_ vssd1 vssd1
+ vccd1 vccd1 _03906_ sky130_fd_sc_hd__or2_1
X_10657_ _06995_ _06996_ _06981_ vssd1 vssd1 vccd1 vccd1 _06997_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_36_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload15 clknet_leaf_158_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload15/Y sky130_fd_sc_hd__inv_16
XFILLER_0_152_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09197__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload26 clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload26/Y sky130_fd_sc_hd__clkinvlp_4
X_16164_ clknet_leaf_134_wb_clk_i net1907 _00152_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13376_ net1581 net829 _03838_ team_01_WB.instance_to_wrap.cpu.f0.i\[1\] vssd1 vssd1
+ vccd1 vccd1 _01871_ sky130_fd_sc_hd__a22o_1
Xclkload37 clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload37/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_77_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09800__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10588_ _06900_ _06910_ vssd1 vssd1 vccd1 vccd1 _06928_ sky130_fd_sc_hd__nor2_4
XFILLER_0_51_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload48 clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload48/Y sky130_fd_sc_hd__clkinv_4
Xclkload59 clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload59/Y sky130_fd_sc_hd__bufinv_16
X_15115_ net1424 vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__inv_2
X_12327_ net3149 net219 net429 vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_149_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16095_ clknet_leaf_126_wb_clk_i _01870_ _00083_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_114_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10961__A2 _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09159__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15046_ net1381 vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__inv_2
X_12258_ _07793_ _07794_ net573 vssd1 vssd1 vccd1 vccd1 _07963_ sky130_fd_sc_hd__and3_1
XFILLER_0_142_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11666__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13854__A_N net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13447__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11209_ net525 _07495_ vssd1 vssd1 vccd1 vccd1 _07549_ sky130_fd_sc_hd__or2_1
XANTENNA__10174__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12189_ net2517 net291 net448 vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__mux2_1
X_16997_ clknet_leaf_52_wb_clk_i _02684_ _00980_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13112__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15948_ net1361 vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__inv_2
XANTENNA__13663__A1 _07639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09660__A net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10477__A1 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09331__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12497__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15879_ net1357 vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__inv_2
X_08420_ net1020 net941 vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__and2_1
X_17618_ clknet_leaf_2_wb_clk_i _03303_ _01559_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_148_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08707__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08351_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[30\] net811 _04642_ _04644_
+ _04689_ vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__a2111o_1
X_17549_ clknet_leaf_68_wb_clk_i _03236_ _01532_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_08282_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[1\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__and2_1
XANTENNA__13179__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload9 clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload9/Y sky130_fd_sc_hd__inv_8
XFILLER_0_116_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_93_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_27_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12926__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09398__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_22_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09538__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14128__C1 _04152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12960__S net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1037_A net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14143__A2 _04254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout497_A net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout202 _07858_ vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13357__A _04483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout213 _07838_ vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__buf_2
Xfanout224 _07827_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10165__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1204_A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout235 net236 vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__clkbuf_2
Xfanout246 _07842_ vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__buf_1
X_09805_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[14\] net785 net770 vssd1
+ vssd1 vccd1 vccd1 _06145_ sky130_fd_sc_hd__a21o_1
Xfanout257 net258 vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input2_A DAT_I[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout268 _07877_ vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__clkbuf_2
Xfanout279 _07917_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__clkbuf_2
X_07997_ team_01_WB.instance_to_wrap.cpu.f0.num\[22\] vssd1 vssd1 vccd1 vccd1 _04495_
+ sky130_fd_sc_hd__inv_2
XANTENNA_fanout664_A _04806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09736_ net996 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[20\] net980 vssd1
+ vssd1 vccd1 vccd1 _06076_ sky130_fd_sc_hd__and3_1
XANTENNA__09858__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13654__A1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09570__A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09322__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09667_ net1136 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[22\] net981
+ vssd1 vssd1 vccd1 vccd1 _06007_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout452_X net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout831_A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14188__A net1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout929_A net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08618_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[11\] net686 net646 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[11\]
+ _04950_ vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__a221o_1
XANTENNA__12200__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13406__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09598_ net1146 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[24\] net985
+ vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__and3_1
XFILLER_0_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11324__B team_01_WB.instance_to_wrap.cpu.DM0.data_i\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08549_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[19\] net693 _04886_ _04887_
+ _04888_ vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout717_X net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11560_ net3094 net1182 net37 vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__a21o_1
XANTENNA__08473__X _04813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10511_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[31\] net772 net739 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06851_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_98_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11491_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[17\] net580 vssd1 vssd1 vccd1
+ vccd1 _07773_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_98_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13230_ net2970 net352 net348 team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1
+ vccd1 vccd1 _01920_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09389__A2 _05726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10442_ net504 _06780_ vssd1 vssd1 vccd1 vccd1 _06782_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12393__A1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08597__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13161_ net1647 net849 net841 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[15\] vssd1
+ vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__a22o_1
XANTENNA__13877__A_N team_01_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10373_ _06710_ _06711_ _06708_ vssd1 vssd1 vccd1 vccd1 _06713_ sky130_fd_sc_hd__o21a_1
X_12112_ net2515 net225 net455 vssd1 vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14134__A2 _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input58_A wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13092_ _03715_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[2\] net853 vssd1 vssd1
+ vccd1 vccd1 _02033_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17735__Q team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12043_ net2940 net259 net465 vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__mux2_1
X_16920_ clknet_leaf_38_wb_clk_i _02607_ _00903_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09464__B _05802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16851_ clknet_leaf_17_wb_clk_i _02538_ _00834_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09183__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout780 net781 vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__buf_6
XFILLER_0_102_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15802_ net1211 vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__inv_2
Xfanout791 net793 vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_4_14__f_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16782_ clknet_leaf_27_wb_clk_i _02469_ _00765_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13645__A1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09849__B1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13994_ _04229_ _04238_ _04247_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[64\]
+ vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_137_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15733_ net1285 vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12945_ net357 _03705_ _03706_ net870 net2281 vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__a32o_1
XFILLER_0_88_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11120__A2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12110__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15664_ net1273 vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__inv_2
X_12876_ net2119 net872 net359 _03658_ vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__a22o_1
X_17403_ clknet_leaf_74_wb_clk_i _03090_ _01386_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08527__C net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14615_ net1337 vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__inv_2
X_11827_ net2039 net189 net487 vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__mux2_1
X_15595_ net1397 vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17334_ clknet_leaf_13_wb_clk_i _03021_ _01317_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11758_ net576 _07794_ _07942_ vssd1 vssd1 vccd1 vccd1 _07943_ sky130_fd_sc_hd__and3_1
X_14546_ net1365 vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10709_ net514 _07024_ _06967_ vssd1 vssd1 vccd1 vccd1 _07049_ sky130_fd_sc_hd__a21boi_1
X_17265_ clknet_leaf_118_wb_clk_i _02952_ _01248_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11689_ net2152 net257 net500 vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_116_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14477_ net1411 vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload104 clknet_leaf_96_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload104/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_102_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16216_ clknet_leaf_139_wb_clk_i net1916 _00204_ vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_144_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13428_ _03887_ _03888_ vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__or2_1
Xclkload115 clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload115/Y sky130_fd_sc_hd__clkinv_2
Xclkload126 clknet_leaf_74_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload126/Y sky130_fd_sc_hd__clkinv_4
X_17196_ clknet_leaf_16_wb_clk_i _02883_ _01179_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload137 clknet_leaf_98_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload137/Y sky130_fd_sc_hd__inv_6
Xclkload148 clknet_leaf_90_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload148/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_51_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08588__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12780__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16147_ clknet_leaf_128_wb_clk_i _01910_ _00135_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13359_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[12\] _03830_ net827 vssd1 vssd1
+ vccd1 vccd1 _01880_ sky130_fd_sc_hd__mux2_1
XANTENNA__10395__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10934__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16078_ clknet_leaf_131_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[0\]
+ _00066_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17645__Q team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15029_ net1276 vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__inv_2
XANTENNA__10147__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09552__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09093__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_140_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_140_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xinput2 DAT_I[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10032__C net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09521_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[29\] net822 net773 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[29\]
+ _05848_ vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__a221o_1
XANTENNA__09304__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09452_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[29\] net685 net678 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[29\]
+ _05785_ vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12020__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08403_ _04732_ _04739_ _04742_ vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__nand3_2
XANTENNA__08437__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10870__A1 _06636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09383_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[26\] net697 net678 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12808__X _03634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout245_A _07842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08334_ net992 net968 vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08265_ net2572 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[8\] net1049 vssd1 vssd1
+ vccd1 vccd1 _03422_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout412_A _03563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1154_A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08196_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[85\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[77\]
+ net1050 vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12690__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08043__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1321_A net1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09565__A net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14116__A2 _04258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08594__A3 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08900__C net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout879_A _04810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11159__X _07499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1008 net1015 vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1019 net1021 vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1207_X net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09543__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout667_X net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08468__X _04808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13627__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09719_ _06055_ _06056_ _06057_ _06058_ vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout834_X net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10991_ net375 _07326_ _07328_ _07330_ _06905_ vssd1 vssd1 vccd1 vccd1 _07331_ sky130_fd_sc_hd__a32o_1
XANTENNA__09731__C net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08503__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11102__A2 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ _04510_ _03579_ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_48_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17001__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12661_ net3111 net208 net389 vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12865__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14400_ net1358 vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_65_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ net1956 net223 net499 vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__mux2_1
X_12592_ net2294 net215 net397 vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__mux2_1
X_15380_ net1380 vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_137_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08644__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14331_ net1326 vssd1 vssd1 vccd1 vccd1 _00125_ sky130_fd_sc_hd__inv_2
X_11543_ net1677 net1173 net590 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\] vssd1
+ vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17050_ clknet_leaf_78_wb_clk_i _02737_ _01033_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_14262_ net1204 vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__inv_2
X_11474_ net366 _07764_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[26\] net874
+ vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_52_269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13213_ net24 net838 net630 net2996 vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__a22o_1
X_16001_ net1410 vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__inv_2
X_10425_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[27\] net801 net754 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06765_ sky130_fd_sc_hd__a22o_1
X_14193_ net3051 _04458_ _04460_ vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__o21a_1
XANTENNA__08034__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_111_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13144_ team_01_WB.instance_to_wrap.a1.curr_state\[1\] _04509_ team_01_WB.instance_to_wrap.a1.curr_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__and3b_4
XANTENNA__09475__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10356_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[17\] net814 _06678_ _06687_
+ _06688_ vssd1 vssd1 vccd1 vccd1 _06696_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09782__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_11__f_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_11__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_13075_ net3084 net3015 net861 vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__mux2_1
X_17952_ net1467 vssd1 vssd1 vccd1 vccd1 gpio_out[35] sky130_fd_sc_hd__buf_2
X_10287_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[19\] net807 net755 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _06627_ sky130_fd_sc_hd__a22o_1
XANTENNA__10414__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12105__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12026_ net2076 net188 net463 vssd1 vssd1 vccd1 vccd1 _02958_ sky130_fd_sc_hd__mux2_1
X_16903_ clknet_leaf_99_wb_clk_i _02590_ _00886_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_17883_ clknet_leaf_139_wb_clk_i _03558_ _01823_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11944__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16834_ clknet_leaf_76_wb_clk_i _02521_ _00817_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13618__A1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_109_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16765_ clknet_leaf_65_wb_clk_i _02452_ _00748_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13977_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[80\] _04251_ _04267_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__a22o_1
X_15716_ net1222 vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12928_ _05490_ _07757_ _03694_ vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__o21ai_1
X_16696_ clknet_leaf_61_wb_clk_i _02383_ _00679_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15647_ net1314 vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__inv_2
X_12859_ net3025 net296 net381 vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__mux2_1
XANTENNA__14043__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08554__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15578_ net1314 vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17317_ clknet_leaf_50_wb_clk_i _03004_ _01300_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_14529_ net1364 vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08050_ team_01_WB.instance_to_wrap.cpu.K0.code\[7\] team_01_WB.instance_to_wrap.cpu.K0.code\[5\]
+ team_01_WB.instance_to_wrap.cpu.K0.code\[4\] team_01_WB.instance_to_wrap.cpu.K0.code\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__or4b_2
X_17248_ clknet_leaf_45_wb_clk_i _02935_ _01231_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09088__C net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17644__CLK clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13554__B1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17179_ clknet_leaf_74_wb_clk_i _02866_ _01162_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10027__C net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09773__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08952_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[6\] net689 _05269_ _05276_
+ _05277_ vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12015__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10324__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11283__D_N _07600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11139__B _06924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08883_ net598 _05219_ _05221_ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout195_A _07634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11854__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_82 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08288__X _04628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13609__A1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout362_A _03580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08448__B net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09504_ net1149 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[29\] net949
+ vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_13__f_wb_clk_i_X clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_78_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09435_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[28\] net696 net663 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__a22o_1
XANTENNA__12685__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1369_A net1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09366_ net598 _05704_ vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_43_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08317_ net1155 net959 vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10058__X _06398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_40 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09297_ net1002 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[22\] net929 vssd1
+ vssd1 vccd1 vccd1 _05637_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout415_X net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_51 _03654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1157_X net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_62 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08248_ net2321 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[25\] net1057 vssd1 vssd1
+ vccd1 vccd1 _03439_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout996_A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08179_ net2872 net2730 net1044 vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10359__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10210_ _06547_ _06548_ _06549_ vssd1 vssd1 vccd1 vccd1 _06550_ sky130_fd_sc_hd__or3_1
XANTENNA__11288__C_N net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09295__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11190_ net328 _07526_ _07529_ net555 _07525_ vssd1 vssd1 vccd1 vccd1 _07530_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout784_X net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10141_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[11\] net815 net779 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06481_ sky130_fd_sc_hd__a22o_1
Xoutput180 net180 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09516__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10072_ net1137 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[7\] net981 vssd1
+ vssd1 vccd1 vccd1 _06412_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout951_X net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08724__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11764__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13900_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[5\] _04201_ vssd1 vssd1 vccd1
+ vccd1 _04202_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_89_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14880_ net1238 vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__inv_2
XANTENNA__08639__A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10531__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13831_ net2026 net831 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[24\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_67_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16550_ clknet_leaf_1_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[16\]
+ _00533_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13762_ _04141_ _04148_ _04149_ _04150_ vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__and4_1
X_10974_ _05301_ net332 _07313_ net336 net369 vssd1 vssd1 vccd1 vccd1 _07314_ sky130_fd_sc_hd__a221o_1
XANTENNA__08926__X _05266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15501_ net1266 vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__inv_2
X_12713_ net2051 net296 net386 vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16481_ clknet_leaf_152_wb_clk_i _02235_ _00464_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12595__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13693_ team_01_WB.instance_to_wrap.cpu.c0.count\[7\] team_01_WB.instance_to_wrap.cpu.c0.count\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__nand2_1
X_15432_ net1376 vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12644_ net3044 net282 net393 vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__mux2_1
XANTENNA__08374__A team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_156_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17667__CLK clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08805__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12575_ net2332 net287 net402 vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15363_ net1249 vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17102_ clknet_leaf_28_wb_clk_i _02789_ _01085_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_152_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14314_ net1325 vssd1 vssd1 vccd1 vccd1 _00108_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_152_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11526_ net1731 net1171 net588 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] vssd1
+ vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__a22o_1
X_15294_ net1320 vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17033_ clknet_leaf_40_wb_clk_i _02720_ _01016_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11939__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11457_ _04712_ _04753_ vssd1 vssd1 vccd1 vccd1 _07753_ sky130_fd_sc_hd__or2_1
X_14245_ net1230 vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10408_ _06598_ _06604_ _06743_ _06107_ vssd1 vssd1 vccd1 vccd1 _06748_ sky130_fd_sc_hd__a211o_1
XFILLER_0_141_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14176_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[9\] _04448_ net1426 vssd1
+ vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_68_48 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11388_ team_01_WB.instance_to_wrap.cpu.f0.i\[30\] _07716_ _07699_ vssd1 vssd1 vccd1
+ vccd1 _07717_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09636__C net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10339_ net1137 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[17\] net963
+ vssd1 vssd1 vccd1 vccd1 _06679_ sky130_fd_sc_hd__and3_1
X_13127_ net1802 net845 net634 team_01_WB.instance_to_wrap.a1.ADR_I\[16\] vssd1 vssd1
+ vccd1 vccd1 _02014_ sky130_fd_sc_hd__a22o_1
X_17935_ team_01_WB.instance_to_wrap.cpu.LCD0.lcd_rs vssd1 vssd1 vccd1 vccd1 net157
+ sky130_fd_sc_hd__clkbuf_1
X_13058_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[28\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[36\]
+ net858 vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_9__f_wb_clk_i_X clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11674__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1350 net1355 vssd1 vssd1 vccd1 vccd1 net1350 sky130_fd_sc_hd__buf_4
X_12009_ net2831 net230 net468 vssd1 vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__mux2_1
Xfanout1361 net1362 vssd1 vssd1 vccd1 vccd1 net1361 sky130_fd_sc_hd__buf_2
X_17866_ clknet_leaf_125_wb_clk_i _03541_ _01806_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_128_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1372 net1373 vssd1 vssd1 vccd1 vccd1 net1372 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_128_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1383 net1384 vssd1 vssd1 vccd1 vccd1 net1383 sky130_fd_sc_hd__buf_4
Xfanout1394 net1398 vssd1 vssd1 vccd1 vccd1 net1394 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16539__Q team_01_WB.instance_to_wrap.cpu.DM0.data_i\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16817_ clknet_leaf_116_wb_clk_i _02504_ _00800_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_17797_ clknet_leaf_95_wb_clk_i net2419 _01737_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[67\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15670__A net1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16748_ clknet_leaf_147_wb_clk_i _02435_ _00731_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_34_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_49_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09691__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[22\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16679_ clknet_leaf_104_wb_clk_i _02366_ _00662_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09220_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[17\] net664 _05533_
+ _05543_ _05549_ vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_29_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08715__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09151_ _05456_ _05490_ net603 vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__mux2_2
XFILLER_0_57_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08102_ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[12\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[15\]
+ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[14\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__or4b_1
XFILLER_0_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09082_ net1011 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[13\] net939 vssd1
+ vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__and3_1
XANTENNA__10053__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire585_X net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09994__A2 _04636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11849__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08033_ net1602 net567 net345 net1069 vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__a22o_1
Xinput60 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_1
Xhold800 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2335 sky130_fd_sc_hd__dlygate4sd3_1
Xinput71 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__buf_1
Xhold811 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[0\] vssd1 vssd1 vccd1 vccd1 net2346
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold822 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2357 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09746__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold833 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold855 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2401 sky130_fd_sc_hd__dlygate4sd3_1
Xhold877 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2412 sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 team_01_WB.instance_to_wrap.cpu.c0.count\[13\] vssd1 vssd1 vccd1 vccd1 net2423
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09984_ _06318_ _06321_ _06322_ _06323_ vssd1 vssd1 vccd1 vccd1 _06324_ sky130_fd_sc_hd__or4_1
Xhold899 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2434 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1117_A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08935_ net1112 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[6\] net894 vssd1
+ vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_73_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout198_X net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1500 team_01_WB.instance_to_wrap.cpu.f0.num\[15\] vssd1 vssd1 vccd1 vccd1 net3035
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout577_A net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11305__A2 _07476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1511 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net3046 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1522 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net3057 sky130_fd_sc_hd__dlygate4sd3_1
X_08866_ net1106 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[3\] net937 vssd1
+ vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__and3_1
Xhold1533 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[40\] vssd1 vssd1 vccd1 vccd1
+ net3068 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1544 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net3079 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1555 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[2\] vssd1 vssd1 vccd1 vccd1
+ net3090 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1566 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[22\] vssd1 vssd1 vccd1 vccd1
+ net3101 sky130_fd_sc_hd__dlygate4sd3_1
X_08797_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[0\] net690 _05134_ _05135_
+ _05136_ vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09281__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1577 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net3112 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1588 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net3123 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout365_X net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1599 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3134 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15580__A net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12805__A2 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10816__A1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout911_A net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout532_X net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14196__A net1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09418_ _05756_ _05757_ net597 vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__mux2_2
XANTENNA__10292__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10690_ net523 _07029_ vssd1 vssd1 vccd1 vccd1 _07030_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12569__A1 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09349_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[25\] net681 net677 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[25\]
+ _05688_ vssd1 vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10044__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11241__A1 _06919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12360_ net2825 net219 net425 vssd1 vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__mux2_1
XANTENNA__09985__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08481__X _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13518__B1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11311_ _04505_ _04524_ vssd1 vssd1 vccd1 vccd1 _07649_ sky130_fd_sc_hd__nor2_1
XANTENNA__11759__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12291_ _07794_ _07942_ net573 vssd1 vssd1 vccd1 vccd1 _07964_ sky130_fd_sc_hd__and3_4
X_14030_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[34\] _04230_ _04236_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[50\]
+ _04311_ vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__a221o_1
X_11242_ _05729_ net330 _07581_ net368 vssd1 vssd1 vccd1 vccd1 _07582_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13259__B net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12741__A1 _07088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11173_ _05417_ net341 net334 _07512_ vssd1 vssd1 vccd1 vccd1 _07513_ sky130_fd_sc_hd__a31o_1
XFILLER_0_140_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10124_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[6\] net765 net624 vssd1
+ vssd1 vccd1 vccd1 _06464_ sky130_fd_sc_hd__o21ai_1
XANTENNA_input40_A wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15981_ net1416 vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__inv_2
X_17720_ clknet_leaf_156_wb_clk_i _00005_ _01661_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10055_ _06391_ _06392_ _06393_ _06394_ vssd1 vssd1 vccd1 vccd1 _06395_ sky130_fd_sc_hd__or4_1
X_14932_ net1379 vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__inv_2
XANTENNA__10504__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09370__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17651_ clknet_leaf_149_wb_clk_i _03336_ _01592_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14863_ net1385 vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__inv_2
XANTENNA__09191__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11507__B _07756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16602_ clknet_leaf_78_wb_clk_i _02289_ _00585_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15490__A net1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13814_ net2158 net832 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[7\]
+ sky130_fd_sc_hd__and2_1
X_17582_ clknet_leaf_96_wb_clk_i _03269_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__dfxtp_1
X_14794_ net1374 vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_123_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16533_ clknet_leaf_157_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[31\]
+ _00516_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13745_ net1181 team_01_WB.instance_to_wrap.cpu.RU0.state\[2\] vssd1 vssd1 vccd1
+ vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_ihit sky130_fd_sc_hd__and2b_1
XFILLER_0_97_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10957_ net335 _06919_ _07296_ vssd1 vssd1 vccd1 vccd1 _07297_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10283__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16464_ clknet_leaf_25_wb_clk_i _02218_ _00447_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13676_ net1688 net569 net347 team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1
+ vccd1 vccd1 _01826_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_118_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10888_ net530 _07227_ _07213_ vssd1 vssd1 vccd1 vccd1 _07228_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15415_ net1221 vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__inv_2
X_12627_ net2991 net245 net392 vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__mux2_1
X_16395_ clknet_leaf_119_wb_clk_i net2961 _00378_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[118\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15346_ net1292 vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__inv_2
X_12558_ net2504 net219 net401 vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__mux2_1
XANTENNA__08832__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13509__B1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10586__A3 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11669__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11509_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[8\] _07756_ vssd1 vssd1 vccd1
+ vccd1 _07782_ sky130_fd_sc_hd__and2_1
X_15277_ net1263 vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__inv_2
Xhold107 _01986_ vssd1 vssd1 vccd1 vccd1 net1642 sky130_fd_sc_hd__dlygate4sd3_1
X_12489_ _07945_ _07951_ net574 vssd1 vssd1 vccd1 vccd1 _03564_ sky130_fd_sc_hd__and3_4
XFILLER_0_80_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold118 net103 vssd1 vssd1 vccd1 vccd1 net1653 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14182__B1 net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17016_ clknet_leaf_27_wb_clk_i _02703_ _00999_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold129 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[25\] vssd1 vssd1 vccd1 vccd1
+ net1664 sky130_fd_sc_hd__dlygate4sd3_1
X_14228_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[4\] vssd1 vssd1 vccd1
+ vccd1 _02259_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11535__A2 net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15665__A net1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14159_ _04187_ _04439_ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout609 _03583_ vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1068 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09663__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08720_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[5\] net682 net678 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_47_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_17918_ net1525 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
Xfanout1180 net1181 vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__buf_2
XANTENNA__09361__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08651_ net1020 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[10\] net919 vssd1
+ vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__and3_1
Xfanout1191 net1192 vssd1 vssd1 vccd1 vccd1 net1191 sky130_fd_sc_hd__buf_2
X_17849_ clknet_leaf_121_wb_clk_i _03525_ _01789_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_157_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08582_ net1104 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[15\] net881
+ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10040__C net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12799__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09203_ net1083 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[17\] net917
+ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout325_A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12816__X _03640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09134_ net1023 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[14\] net931 vssd1
+ vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1067_A team_01_WB.instance_to_wrap.cpu.RU0.state\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09967__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11223__B2 _05263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11579__S net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09065_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[12\] net666 _05388_
+ _05396_ _05404_ vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08461__B net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1234_A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08016_ team_01_WB.instance_to_wrap.cpu.K0.code\[6\] team_01_WB.instance_to_wrap.cpu.K0.code\[5\]
+ team_01_WB.instance_to_wrap.cpu.K0.code\[4\] team_01_WB.instance_to_wrap.cpu.K0.code\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__or4b_2
Xhold630 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2165 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout694_A net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold641 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2176 sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2187 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold663 _01991_ vssd1 vssd1 vccd1 vccd1 net2198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2220 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1022_X net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold696 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2231 sky130_fd_sc_hd__dlygate4sd3_1
X_09967_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[3\] net809 net732 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06307_ sky130_fd_sc_hd__a22o_1
XANTENNA__13807__B net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout861_A net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout482_X net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11167__X _07507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout959_A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08918_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[2\] net704 _05253_ _05257_
+ vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__o22a_4
XANTENNA__12203__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09898_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[5\] net731 _06222_ _06226_
+ _06230_ vssd1 vssd1 vccd1 vccd1 _06238_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_86_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1330 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2865 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09352__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1341 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[88\] vssd1 vssd1 vccd1 vccd1
+ net2876 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1352 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2887 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1363 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[98\] vssd1 vssd1 vccd1 vccd1
+ net2898 sky130_fd_sc_hd__dlygate4sd3_1
X_08849_ net599 _05187_ _05188_ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout747_X net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1374 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2909 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1385 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2920 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1396 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2931 sky130_fd_sc_hd__dlygate4sd3_1
X_11860_ net2186 net190 net483 vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10811_ _06969_ _07150_ _07140_ vssd1 vssd1 vccd1 vccd1 _07151_ sky130_fd_sc_hd__o21ai_2
XANTENNA__13987__B1 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11791_ _07790_ net575 _07794_ vssd1 vssd1 vccd1 vccd1 _07944_ sky130_fd_sc_hd__and3_4
XANTENNA__09655__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[23\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout914_X net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11343__A team_01_WB.instance_to_wrap.cpu.f0.i\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13530_ net721 _07579_ net1074 vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__o21a_1
XANTENNA__11462__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10742_ _07080_ _07081_ net515 vssd1 vssd1 vccd1 vccd1 _07082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13461_ _03854_ _03855_ vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__nor2_1
X_10673_ net552 _06340_ _07012_ vssd1 vssd1 vccd1 vccd1 _07013_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08923__Y _05263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11630__X _07842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15200_ net1235 vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12412_ net2551 net249 net422 vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__mux2_1
XANTENNA__10017__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09958__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16180_ clknet_leaf_7_wb_clk_i _01940_ _00168_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08652__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13392_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] _04885_ vssd1 vssd1
+ vccd1 vccd1 _03853_ sky130_fd_sc_hd__or2_1
XFILLER_0_152_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15131_ net1253 vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__inv_2
XANTENNA__12962__A1 _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12343_ net1931 net254 net428 vssd1 vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08091__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15062_ net1258 vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__inv_2
X_12274_ net2971 net263 net436 vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14013_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[41\] _04256_ _04263_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[121\]
+ _04291_ vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__a221o_1
X_11225_ _06934_ _07201_ _07562_ _07564_ vssd1 vssd1 vccd1 vccd1 _07565_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_75_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11156_ net530 _07495_ vssd1 vssd1 vccd1 vccd1 _07496_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_147_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10107_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[6\] net781 net741 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06447_ sky130_fd_sc_hd__a22o_1
XANTENNA__12113__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11087_ _05781_ _05899_ _07045_ _07426_ vssd1 vssd1 vccd1 vccd1 _07427_ sky130_fd_sc_hd__a31o_1
X_15964_ net1366 vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__inv_2
XANTENNA__10422__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_125_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17703_ clknet_leaf_134_wb_clk_i _03387_ _01644_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[24\]
+ sky130_fd_sc_hd__dfrtp_4
X_10038_ net1142 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[0\] net958 vssd1
+ vssd1 vccd1 vccd1 _06378_ sky130_fd_sc_hd__and3_1
X_14915_ net1250 vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__inv_2
XANTENNA__08697__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15895_ net1413 vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__inv_2
XANTENNA__11952__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17634_ clknet_leaf_157_wb_clk_i _03319_ _01575_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_19_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14846_ net1345 vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_121_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08827__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13978__B1 _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17565_ clknet_leaf_88_wb_clk_i _03252_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14777_ net1237 vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__inv_2
X_11989_ net2074 net318 net474 vssd1 vssd1 vccd1 vccd1 _02993_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16516_ clknet_leaf_1_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[14\]
+ _00499_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13728_ net1170 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[4\] team_01_WB.instance_to_wrap.cpu.DM0.enable
+ _04711_ vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__or4_1
XANTENNA__11453__A1 net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17496_ clknet_leaf_50_wb_clk_i _03183_ _01479_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16447_ clknet_leaf_78_wb_clk_i _02201_ _00430_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12783__S net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13659_ net727 net321 net988 vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_140_Right_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11205__A1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10008__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09658__A _04844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16378_ clknet_leaf_101_wb_clk_i _02132_ _00361_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[101\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_30_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08082__A0 team_01_WB.instance_to_wrap.cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_124_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11700__B net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15329_ net1280 vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__inv_2
XANTENNA__17385__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10964__B1 _07300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09096__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11508__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10035__C net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout406 _03565_ vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__buf_6
X_09821_ _05491_ _06160_ vssd1 vssd1 vccd1 vccd1 _06161_ sky130_fd_sc_hd__xor2_1
XANTENNA__09582__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout417 _03562_ vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__clkbuf_8
Xfanout428 _07965_ vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__buf_4
Xfanout439 _07962_ vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12023__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09752_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[20\] net805 net737 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__a22o_1
XANTENNA__10332__A _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08703_ net602 net585 _05041_ vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__a21oi_2
X_09683_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[22\] net801 net799 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06023_ sky130_fd_sc_hd__a22o_1
XANTENNA__12958__S net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout275_A _07851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11862__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08634_ net1020 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[10\] net908
+ vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__and3_1
XANTENNA__08296__X _04636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08737__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08565_ net999 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[19\] net944 vssd1
+ vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout442_A _07962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1184_A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10247__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08496_ _04827_ _04828_ _04829_ _04835_ vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__or4_2
XFILLER_0_76_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10798__A3 _06811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12693__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1351_A net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout707_A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout328_X net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08903__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09117_ net1110 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[14\] net898
+ vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__and3_1
XANTENNA__08073__B1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08612__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09048_ net1029 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[12\] net885 vssd1
+ vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout697_X net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold460 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[6\] vssd1 vssd1 vccd1 vccd1
+ net1995 sky130_fd_sc_hd__dlygate4sd3_1
Xhold471 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[8\] vssd1 vssd1 vccd1 vccd1
+ net2006 sky130_fd_sc_hd__dlygate4sd3_1
Xhold482 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2017 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ _05682_ net511 vssd1 vssd1 vccd1 vccd1 _07350_ sky130_fd_sc_hd__nor2_1
XANTENNA__08376__A1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold493 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2028 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09734__C net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout940 _04759_ vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__buf_4
Xfanout951 _04662_ vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout973 net974 vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__clkbuf_2
Xfanout984 _04629_ vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout995 _04491_ vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09325__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12961_ net1938 net870 net357 _03715_ vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_142_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09876__A1 _06215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1160 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2695 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13672__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11772__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1171 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2706 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11625__X _07838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14700_ net1210 vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__inv_2
X_11912_ net3031 net286 net482 vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__mux2_1
Xhold1182 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2717 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11683__A1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15680_ net1242 vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__inv_2
XANTENNA__08647__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1193 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2728 sky130_fd_sc_hd__dlygate4sd3_1
X_12892_ _05678_ net577 vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__nor2_1
X_14631_ net1374 vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11843_ net3024 net231 net489 vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11073__A _05566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10238__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17350_ clknet_leaf_72_wb_clk_i _03037_ _01333_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14562_ net1366 vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__inv_2
X_11774_ net2211 net264 net498 vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16301_ clknet_leaf_123_wb_clk_i _02055_ _00284_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13513_ net721 _07088_ net1074 vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__o21a_1
XFILLER_0_27_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17281_ clknet_leaf_54_wb_clk_i _02968_ _01264_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10725_ _07060_ _07064_ net529 vssd1 vssd1 vccd1 vccd1 _07065_ sky130_fd_sc_hd__mux2_1
XANTENNA__12456__X _03563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14493_ net1411 vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16232_ clknet_leaf_135_wb_clk_i net1610 _00220_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__dfrtp_1
X_13444_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] _05419_ vssd1 vssd1
+ vccd1 vccd1 _03905_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10656_ net523 _06988_ _06991_ _06906_ net338 vssd1 vssd1 vccd1 vccd1 _06996_ sky130_fd_sc_hd__o221a_1
XFILLER_0_152_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11738__A2 _07449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16163_ clknet_leaf_134_wb_clk_i _01926_ _00151_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[26\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload16 clknet_leaf_159_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload16/Y sky130_fd_sc_hd__inv_6
XANTENNA__11520__B net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10587_ _06883_ net336 _06916_ _06926_ vssd1 vssd1 vccd1 vccd1 _06927_ sky130_fd_sc_hd__a211o_1
XFILLER_0_35_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13375_ net1582 net829 _03838_ team_01_WB.instance_to_wrap.cpu.f0.i\[2\] vssd1 vssd1
+ vccd1 vccd1 _01872_ sky130_fd_sc_hd__a22o_1
Xclkload27 clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload27/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_77_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12108__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload38 clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload38/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_77_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10417__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload49 clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload49/Y sky130_fd_sc_hd__clkinv_4
X_15114_ net1374 vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12326_ net2649 net221 net427 vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_149_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16094_ clknet_leaf_131_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[16\]
+ _00082_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[16\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_114_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11947__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15045_ net1288 vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_114_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12257_ net2635 net290 net440 vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11208_ _06920_ _07050_ _07026_ vssd1 vssd1 vccd1 vccd1 _07548_ sky130_fd_sc_hd__a21bo_1
XANTENNA__13447__B _05380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12188_ net2031 net316 net449 vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__mux2_1
X_11139_ net516 _06924_ vssd1 vssd1 vccd1 vccd1 _07479_ sky130_fd_sc_hd__nor2_1
X_16996_ clknet_leaf_83_wb_clk_i _02683_ _00979_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13648__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09316__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09941__A _06280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15947_ net1367 vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__inv_2
XANTENNA__13463__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15878_ net1348 vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__inv_2
X_14829_ net1265 vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__inv_2
X_17617_ clknet_leaf_2_wb_clk_i _03302_ _01558_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10229__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08350_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[30\] net799 net777 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__a22o_1
X_17548_ clknet_leaf_147_wb_clk_i _03235_ _01531_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08281_ net2346 net1985 net1046 vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__mux2_1
X_17479_ clknet_leaf_107_wb_clk_i _03166_ _01462_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12807__A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09388__A net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_4_Left_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08723__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16282__Q team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12018__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14128__B1 _04396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11857__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_62_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09555__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout203 _07855_ vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__buf_2
Xfanout214 net217 vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__buf_2
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout392_A net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout225 net228 vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__buf_2
Xfanout236 _07873_ vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__clkbuf_2
X_09804_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[14\] net805 net795 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06144_ sky130_fd_sc_hd__a22o_1
Xfanout247 _07842_ vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__buf_2
Xfanout258 _07888_ vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__clkbuf_2
Xfanout269 _07866_ vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__buf_2
X_07996_ team_01_WB.instance_to_wrap.cpu.f0.num\[28\] vssd1 vssd1 vccd1 vccd1 _04494_
+ sky130_fd_sc_hd__inv_2
X_09735_ net1145 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[20\] net952
+ vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__and3_1
XANTENNA__12688__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout657_A _04815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13654__A2 _07449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1399_A net1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10468__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09666_ net1136 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[22\] net954
+ vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__and3_1
XANTENNA__08467__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10297__B1_N _04919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08617_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[11\] net695 net664 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[11\]
+ _04956_ vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__a221o_1
XANTENNA__13406__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09597_ net1145 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[24\] net971
+ vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout445_X net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11324__C team_01_WB.instance_to_wrap.cpu.DM0.data_i\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08548_ net1077 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[19\] net925
+ vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__and3_1
XFILLER_0_65_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout612_X net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13820__B net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08479_ net1112 net898 vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__and2_2
XFILLER_0_9_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11180__X _07520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10510_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[31\] net821 _06830_ _06833_
+ _06841_ vssd1 vssd1 vccd1 vccd1 _06850_ sky130_fd_sc_hd__a2111o_1
X_11490_ net366 _07772_ net3117 net875 vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_98_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08633__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10441_ net504 _06780_ vssd1 vssd1 vccd1 vccd1 _06781_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_21_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13590__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14119__B1 _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10372_ _06708_ _06710_ _06711_ vssd1 vssd1 vccd1 vccd1 _06712_ sky130_fd_sc_hd__or3_1
X_13160_ net115 net847 net839 net1579 vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout981_X net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12111_ net1969 net284 net457 vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__mux2_1
XANTENNA__11767__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_10__f_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_10__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_13091_ _03714_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[3\] net852 vssd1 vssd1
+ vccd1 vccd1 _02034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_72_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09546__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12042_ net3047 net232 net465 vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__mux2_1
Xhold290 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1825 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_144_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16850_ clknet_leaf_110_wb_clk_i _02537_ _00833_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout770 _04672_ vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__clkbuf_8
X_15801_ net1217 vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__inv_2
Xfanout781 _04663_ vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__buf_4
Xfanout792 net793 vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__clkbuf_8
X_16781_ clknet_leaf_109_wb_clk_i _02468_ _00764_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12598__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09849__A1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13993_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[88\] _04240_ _04243_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[24\]
+ _04284_ vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__a221o_1
XANTENNA__13645__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15732_ net1384 vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__inv_2
X_12944_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[9\] net1039 vssd1 vssd1 vccd1
+ vccd1 _03706_ sky130_fd_sc_hd__or2_1
XANTENNA__10459__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15663_ net1388 vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__inv_2
X_12875_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[30\] _03657_ net1040 vssd1
+ vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__mux2_1
X_17402_ clknet_leaf_79_wb_clk_i _03089_ _01385_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11408__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14614_ net1310 vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__inv_2
X_11826_ net575 _07945_ _07946_ vssd1 vssd1 vccd1 vccd1 _07947_ sky130_fd_sc_hd__and3_4
X_15594_ net1283 vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__inv_2
XANTENNA__14070__A2 _04226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17333_ clknet_leaf_118_wb_clk_i _03020_ _01316_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14545_ net1411 vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__inv_2
X_11757_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\] team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\]
+ vssd1 vssd1 vccd1 vccd1 _07942_ sky130_fd_sc_hd__and2b_2
XFILLER_0_71_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10092__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10708_ _06912_ _07045_ _07047_ vssd1 vssd1 vccd1 vccd1 _07048_ sky130_fd_sc_hd__o21ai_1
X_17264_ clknet_leaf_146_wb_clk_i _02951_ _01247_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14476_ net1416 vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11688_ net612 _07810_ _07887_ _07886_ vssd1 vssd1 vccd1 vccd1 _07888_ sky130_fd_sc_hd__a31o_4
XANTENNA__09639__C net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12908__A1 _03680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16215_ clknet_leaf_124_wb_clk_i net1900 _00203_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__dfrtp_1
X_13427_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] _04971_ vssd1 vssd1
+ vccd1 vccd1 _03888_ sky130_fd_sc_hd__xor2_1
Xclkload105 clknet_leaf_97_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload105/Y sky130_fd_sc_hd__inv_8
Xclkload116 clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload116/X sky130_fd_sc_hd__clkbuf_8
X_10639_ net523 _06928_ vssd1 vssd1 vccd1 vccd1 _06979_ sky130_fd_sc_hd__and2_1
X_17195_ clknet_leaf_9_wb_clk_i _02882_ _01178_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload127 clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload127/Y sky130_fd_sc_hd__inv_6
XFILLER_0_144_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13581__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09495__X _05835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload138 clknet_leaf_100_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload138/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16146_ clknet_leaf_128_wb_clk_i _01909_ _00134_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13358_ net586 _07686_ _03829_ _03828_ net565 vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__a32o_1
XFILLER_0_122_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12309_ net2306 net260 net433 vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16077_ clknet_leaf_130_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_atmax _00065_
+ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.enable sky130_fd_sc_hd__dfrtp_1
X_13289_ team_01_WB.instance_to_wrap.cpu.f0.i\[24\] _03751_ vssd1 vssd1 vccd1 vccd1
+ _03776_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15028_ net1378 vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11895__A1 _07831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09671__A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput3 DAT_I[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
X_16979_ clknet_leaf_24_wb_clk_i _02666_ _00962_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_09520_ _05856_ _05857_ _05858_ _05859_ vssd1 vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__or4_1
XFILLER_0_127_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12301__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08718__C net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09451_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[29\] net669 _05782_ _05789_
+ _05790_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_148_214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08402_ net1169 _04727_ vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__nand2_1
XANTENNA__10870__A2 _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09382_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[26\] net943 net663 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[26\]
+ net706 vssd1 vssd1 vccd1 vccd1 _05722_ sky130_fd_sc_hd__a221o_1
XANTENNA__09068__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14061__A2 _04246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08276__A0 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08333_ net998 net946 vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__nand2_1
XANTENNA__12072__A1 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_49_Left_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10083__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08264_ net2429 net2328 net1056 vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09225__C1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08195_ net2746 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[78\] net1044 vssd1 vssd1
+ vccd1 vccd1 _03492_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12824__X _03646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout405_A net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08579__A1 _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1147_A net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09776__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08750__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09240__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09284__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_58_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1009 net1010 vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout395_X net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1102_X net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13815__B net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout941_A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout562_X net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07979_ team_01_WB.instance_to_wrap.cpu.f0.i\[17\] vssd1 vssd1 vccd1 vccd1 _04477_
+ sky130_fd_sc_hd__inv_2
X_09718_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[21\] net740 _06037_ _06045_
+ _06047_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12907__B1_N net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12211__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10990_ _07318_ _07329_ net540 vssd1 vssd1 vccd1 vccd1 _07330_ sky130_fd_sc_hd__mux2_1
XANTENNA__08503__A1 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09649_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[23\] net734 _05976_ _05978_
+ _05979_ vssd1 vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__a2111o_1
XANTENNA__14037__C1 _04152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12660_ net3078 net245 net389 vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_67_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _07824_ _07826_ net611 vssd1 vssd1 vccd1 vccd1 _07827_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12591_ net3060 net219 net397 vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13042__S net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14330_ net1202 vssd1 vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11542_ net1805 team_01_WB.instance_to_wrap.cpu.DM0.ihit _07785_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_924 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14261_ net1202 vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__inv_2
X_11473_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[26\] net579 vssd1 vssd1 vccd1
+ vccd1 _07764_ sky130_fd_sc_hd__nand2_1
XANTENNA__12881__S net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16000_ net1411 vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__inv_2
XANTENNA_input70_A wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13212_ net27 net838 net630 net2664 vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__a22o_1
XANTENNA__09756__A net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10424_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[27\] net794 _06751_ _06756_
+ _06758_ vssd1 vssd1 vccd1 vccd1 _06764_ sky130_fd_sc_hd__a2111o_1
X_14192_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[15\] _04458_ net1427 vssd1
+ vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13143_ net75 net844 net632 net1620 vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__a22o_1
X_10355_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[17\] net782 _06681_ _06682_
+ _06686_ vssd1 vssd1 vccd1 vccd1 _06695_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_111_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_76_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09519__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17951_ net1466 vssd1 vssd1 vccd1 vccd1 gpio_out[34] sky130_fd_sc_hd__buf_2
X_10286_ _06622_ _06623_ _06624_ _06625_ vssd1 vssd1 vccd1 vccd1 _06626_ sky130_fd_sc_hd__or4_1
X_13074_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[12\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[20\]
+ net854 vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__mux2_1
XANTENNA__09194__C net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16902_ clknet_leaf_90_wb_clk_i _02589_ _00885_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12025_ net576 _07942_ _07951_ vssd1 vssd1 vccd1 vccd1 _07954_ sky130_fd_sc_hd__and3_4
X_17882_ clknet_leaf_133_wb_clk_i _03557_ _01822_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10133__C net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16833_ clknet_leaf_53_wb_clk_i _02520_ _00816_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09922__C net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12121__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16764_ clknet_leaf_60_wb_clk_i _02451_ _00747_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_109_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13976_ _04219_ _04220_ _04237_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__and3_4
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_24_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15715_ net1252 vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__inv_2
X_12927_ net1041 _03652_ vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__and2_2
X_16695_ clknet_leaf_14_wb_clk_i _02382_ _00678_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_85_Left_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11960__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11061__A2_N _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15646_ net1350 vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__inv_2
X_12858_ net1832 net278 net379 vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__mux2_1
XANTENNA__14043__A2 _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11809_ net2625 net257 net493 vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15577_ net1240 vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__inv_2
X_12789_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[13\] _07553_ net1033 vssd1 vssd1
+ vccd1 vccd1 _03621_ sky130_fd_sc_hd__mux2_1
X_17316_ clknet_leaf_82_wb_clk_i _03003_ _01299_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11801__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14528_ net1352 vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17247_ clknet_leaf_43_wb_clk_i _02934_ _01230_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14459_ net1227 vssd1 vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13554__A1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09758__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10308__C net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17178_ clknet_leaf_78_wb_clk_i _02865_ _01161_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xmax_cap712 _04726_ vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__buf_1
XANTENNA__09222__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_94_Left_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16129_ clknet_leaf_127_wb_clk_i _00020_ _00117_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13306__A1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08951_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[6\] net653 _05279_ _05281_
+ _05284_ vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__a2111o_1
XANTENNA_clkbuf_leaf_63_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_138_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08882_ net598 _05219_ _05221_ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09930__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13609__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12031__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08448__C net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09503_ net997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[29\] net959 vssd1
+ vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__and3_1
XANTENNA__14019__C1 net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13867__A_N net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12819__X _03642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11870__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1097_A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09434_ _05767_ _05769_ _05771_ _05773_ vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__or4_1
XANTENNA__08745__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14034__A2 _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09365_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\] net710 _04841_ vssd1 vssd1
+ vccd1 vccd1 _05705_ sky130_fd_sc_hd__a21o_2
XANTENNA_fanout522_A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1264_A net1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08464__B net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08316_ net1158 net1161 net1166 net1164 vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__nor4b_2
XFILLER_0_19_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_30 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_7_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09296_ net1083 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[22\] net929
+ vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__and3_1
XFILLER_0_145_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_41 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09461__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_52 _03654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_941 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_63 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08247_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[34\] net2212 net1052 vssd1 vssd1
+ vccd1 vccd1 _03440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout408_X net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08178_ net2824 net2640 net1047 vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout891_A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08957__D1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12206__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10140_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[11\] net776 net745 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[11\]
+ _06479_ vssd1 vssd1 vccd1 vccd1 _06480_ sky130_fd_sc_hd__a221o_1
Xoutput170 net170 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__clkbuf_4
Xoutput181 net181 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout777_X net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10071_ net1138 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[7\] net950 vssd1
+ vssd1 vccd1 vccd1 _06411_ sky130_fd_sc_hd__and3_1
XANTENNA__08479__X _04819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09921__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout944_X net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09742__C net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13830_ net2241 net830 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[23\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__11346__A team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13761_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[7\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[6\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[9\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__and4bb_1
X_10973_ _05301_ net372 vssd1 vssd1 vccd1 vccd1 _07313_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11780__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15500_ net1259 vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__inv_2
X_12712_ net1873 net276 net384 vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__mux2_1
X_16480_ clknet_leaf_152_wb_clk_i _02234_ _00463_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13692_ _04112_ _04113_ _04114_ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__or3_1
XANTENNA__14025__A2 _04226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_108_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15431_ net1389 vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__inv_2
X_12643_ net2543 net250 net393 vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_156_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10249__X _06589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_156_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08374__B net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09988__B1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11244__C1 _06903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15362_ net1319 vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__inv_2
X_12574_ net2406 net254 net400 vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09452__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17101_ clknet_leaf_109_wb_clk_i _02788_ _01084_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_14313_ net1325 vssd1 vssd1 vccd1 vccd1 _00107_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_152_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11525_ net1841 net1171 net588 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\] vssd1
+ vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__a22o_1
X_15293_ net1241 vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13536__A1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17032_ clknet_leaf_66_wb_clk_i _02719_ _01015_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input73_X net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14244_ net1236 vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11456_ _04712_ _04753_ vssd1 vssd1 vccd1 vccd1 _07752_ sky130_fd_sc_hd__nor2_4
XANTENNA__08390__A _04708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08821__C net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10407_ _06641_ _06677_ _06745_ _06746_ _06639_ vssd1 vssd1 vccd1 vccd1 _06747_ sky130_fd_sc_hd__o311a_1
XANTENNA__12116__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14175_ _04448_ _04449_ vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11387_ _04466_ _07715_ vssd1 vssd1 vccd1 vccd1 _07716_ sky130_fd_sc_hd__nor2_1
X_13126_ net83 net843 net631 net1545 vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__a22o_1
X_10338_ net993 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[17\] net984 vssd1
+ vssd1 vccd1 vccd1 _06678_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_119_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_119_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11955__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17934_ team_01_WB.instance_to_wrap.cpu.LCD0.lcd_en vssd1 vssd1 vccd1 vccd1 net156
+ sky130_fd_sc_hd__clkbuf_1
X_13057_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[29\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[37\]
+ net859 vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__mux2_1
X_10269_ net1128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[19\] net954
+ vssd1 vssd1 vccd1 vccd1 _06609_ sky130_fd_sc_hd__and3_1
XFILLER_0_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1340 net1343 vssd1 vssd1 vccd1 vccd1 net1340 sky130_fd_sc_hd__buf_4
X_12008_ net2362 net263 net468 vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__mux2_1
XANTENNA__09912__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1351 net1355 vssd1 vssd1 vccd1 vccd1 net1351 sky130_fd_sc_hd__buf_4
X_17865_ clknet_leaf_125_wb_clk_i _03540_ _01805_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1362 net1369 vssd1 vssd1 vccd1 vccd1 net1362 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_128_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1373 net1429 vssd1 vssd1 vccd1 vccd1 net1373 sky130_fd_sc_hd__buf_2
Xfanout1384 net1429 vssd1 vssd1 vccd1 vccd1 net1384 sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_147_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1395 net1397 vssd1 vssd1 vccd1 vccd1 net1395 sky130_fd_sc_hd__buf_4
X_16816_ clknet_leaf_20_wb_clk_i _02503_ _00799_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10160__A net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17796_ clknet_leaf_91_wb_clk_i net2433 _01736_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12786__S net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16747_ clknet_leaf_5_wb_clk_i _02434_ _00730_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13959_ _04219_ _04227_ _04237_ vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__and3_4
XANTENNA__11690__S net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16678_ clknet_leaf_91_wb_clk_i _02365_ _00661_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14016__A2 _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15629_ net1268 vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09979__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13775__A1 team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09150_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[14\] net703 _05486_ _05489_
+ vssd1 vssd1 vccd1 vccd1 _05490_ sky130_fd_sc_hd__o22ai_4
XANTENNA__09099__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08101_ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[9\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[8\]
+ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[11\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__or4_1
XANTENNA__08377__C_N team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09081_ net1012 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[13\] net901
+ vssd1 vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12815__A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10038__C net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08032_ net1855 net567 net345 team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1
+ vccd1 vccd1 _03559_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput50 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_1
Xinput61 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__buf_1
Xinput72 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__buf_1
XANTENNA__11538__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold801 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[75\] vssd1 vssd1 vccd1 vccd1
+ net2336 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold812 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold823 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2358 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold834 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2369 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12026__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold845 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2391 sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2402 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold878 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2413 sky130_fd_sc_hd__dlygate4sd3_1
X_09983_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[2\] net823 net800 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06323_ sky130_fd_sc_hd__a22o_1
Xhold889 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2424 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11865__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11718__X _07912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08934_ net1027 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[6\] net907 vssd1
+ vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1012_A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09903__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1501 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net3036 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1512 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net3047 sky130_fd_sc_hd__dlygate4sd3_1
X_08865_ net1106 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[3\] net894 vssd1
+ vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout472_A _07952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1523 team_01_WB.instance_to_wrap.cpu.f0.num\[10\] vssd1 vssd1 vccd1 vccd1 net3058
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1534 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[8\] vssd1 vssd1 vccd1 vccd1
+ net3069 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1545 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net3080 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1556 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net3091 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1567 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net3102 sky130_fd_sc_hd__dlygate4sd3_1
X_08796_ net1009 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[0\] net934 vssd1
+ vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_28_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1578 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net3113 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_28_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10501__C net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1589 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net3124 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12696__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_154_Right_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout737_A net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1381_A net1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout358_X net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13381__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10816__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08475__A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14007__A2 _04230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09682__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08906__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09417_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] net710 net594 vssd1 vssd1
+ vccd1 vccd1 _05757_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_62_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout904_A _04785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11105__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09348_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[25\] net697 net694 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09279_ _05618_ vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_130_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13518__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11310_ _07648_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] _07638_ vssd1
+ vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12290_ net1955 net288 net436 vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout894_X net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09737__C net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08641__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11241_ net335 _06919_ _07346_ vssd1 vssd1 vccd1 vccd1 _07581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11172_ _05417_ net341 net335 vssd1 vssd1 vccd1 vccd1 _07512_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11775__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10123_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[6\] net810 _06457_ _06461_
+ _06462_ vssd1 vssd1 vccd1 vccd1 _06463_ sky130_fd_sc_hd__a2111oi_2
X_15980_ net1368 vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14931_ net1392 vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__inv_2
X_10054_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[0\] net742 _06374_ _06375_
+ _06378_ vssd1 vssd1 vccd1 vccd1 _06394_ sky130_fd_sc_hd__a2111o_1
XANTENNA_input33_A DAT_I[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09472__C net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11701__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08369__B net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14862_ net1299 vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17650_ clknet_leaf_150_wb_clk_i _03335_ _01591_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10411__C net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16601_ clknet_leaf_104_wb_clk_i _02288_ _00584_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13813_ net1601 net833 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[6\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__17634__CLK clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17581_ clknet_leaf_121_wb_clk_i _03268_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__dfxtp_1
X_14793_ net1293 vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16532_ clknet_leaf_159_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[30\]
+ _00515_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_123_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13744_ team_01_WB.instance_to_wrap.cpu.RU0.state\[6\] net1065 net1181 vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_dhit sky130_fd_sc_hd__o21ba_1
X_10956_ _05043_ _06438_ vssd1 vssd1 vccd1 vccd1 _07296_ sky130_fd_sc_hd__and2_1
XANTENNA__08385__A team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08816__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16463_ clknet_leaf_110_wb_clk_i _02217_ _00446_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13675_ net1681 net567 net345 team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1
+ vccd1 vccd1 _01827_ sky130_fd_sc_hd__a22o_1
X_10887_ net514 _07023_ _07215_ vssd1 vssd1 vccd1 vccd1 _07227_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_14_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15414_ net1255 vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__inv_2
X_12626_ net2829 net211 net391 vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16394_ clknet_leaf_101_wb_clk_i _02148_ _00377_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[117\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__09425__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15345_ net1422 vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12557_ net2901 net223 net399 vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15011__A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13509__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11508_ net1720 net877 _07758_ _07781_ vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__o22a_1
XFILLER_0_80_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15276_ net1257 vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__inv_2
X_12488_ net2959 net291 net412 vssd1 vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__mux2_1
Xhold108 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 net1643
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10991__A1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09189__A1 _05528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17015_ clknet_leaf_14_wb_clk_i _02702_ _00998_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08551__C net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold119 _02004_ vssd1 vssd1 vccd1 vccd1 net1654 sky130_fd_sc_hd__dlygate4sd3_1
X_14227_ net3041 vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__clkbuf_1
X_11439_ net1072 _07676_ vssd1 vssd1 vccd1 vccd1 _07744_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12732__A2 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09944__A _06280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14158_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[1\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[0\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[2\] vssd1 vssd1 vccd1 vccd1 _04439_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13109_ team_01_WB.instance_to_wrap.a1.curr_state\[2\] team_01_WB.instance_to_wrap.a1.curr_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__nor2_1
X_14089_ net3107 net604 vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_76 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17917_ net1524 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
XANTENNA__10602__B _06526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1170 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[6\] vssd1 vssd1 vccd1 vccd1
+ net1170 sky130_fd_sc_hd__buf_2
X_08650_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[10\] net932
+ vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__and3_1
Xfanout1181 team_01_WB.instance_to_wrap.a1.BUSY_O vssd1 vssd1 vccd1 vccd1 net1181
+ sky130_fd_sc_hd__clkbuf_2
Xfanout1192 net1207 vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__buf_2
X_17848_ clknet_leaf_119_wb_clk_i net2455 _01788_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[118\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08847__X _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10321__C net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08581_ net1104 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[15\] net895
+ vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_87_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_17779_ clknet_leaf_94_wb_clk_i net2382 _01719_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09113__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[13\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12799__A2 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_16_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09202_ net1085 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[17\] net944
+ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_22_Left_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09416__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09133_ net1022 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[14\] net893
+ vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11223__A2 _06906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08624__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout220_A _07831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10431__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09064_ net1113 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[12\] net899
+ vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10982__A1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10982__B2 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08015_ _04504_ team_01_WB.instance_to_wrap.cpu.f0.state\[7\] vssd1 vssd1 vccd1 vccd1
+ _04511_ sky130_fd_sc_hd__and2_1
Xhold620 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold642 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2177 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1227_A net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold653 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2188 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold664 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2199 sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2210 sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2221 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold697 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2232 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout687_A _04776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09966_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[3\] net796 _06288_ _06289_
+ _06294_ vssd1 vssd1 vccd1 vccd1 _06306_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_31_Left_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1015_X net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08917_ _05248_ _05254_ _05255_ _05256_ vssd1 vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__or4_1
XANTENNA__09292__C net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09897_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[5\] net735 _06225_ _06228_
+ _06229_ vssd1 vssd1 vccd1 vccd1 _06237_ sky130_fd_sc_hd__a2111o_1
Xhold1320 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2855 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout475_X net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1331 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2866 sky130_fd_sc_hd__dlygate4sd3_1
X_08848_ net601 _05153_ _05154_ vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_51_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1342 _03494_ vssd1 vssd1 vccd1 vccd1 net2877 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1353 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2888 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1364 _02129_ vssd1 vssd1 vccd1 vccd1 net2899 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1375 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[91\] vssd1 vssd1 vccd1 vccd1
+ net2910 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1386 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[9\] vssd1 vssd1 vccd1 vccd1
+ net2921 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13823__B net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08779_ net1009 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[0\] net905 vssd1
+ vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__and3_1
Xhold1397 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2932 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1384_X net1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ net529 net516 vssd1 vssd1 vccd1 vccd1 _07150_ sky130_fd_sc_hd__nand2_1
X_11790_ net2293 net290 net498 vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08636__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10741_ _06983_ _06985_ net536 vssd1 vssd1 vccd1 vccd1 _07081_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_40_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11462__A2 _07757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout907_X net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13460_ _03856_ _03858_ _03919_ _04847_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\]
+ vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__a32o_1
X_10672_ net552 _06366_ vssd1 vssd1 vccd1 vccd1 _07012_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09407__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12411_ net2708 net227 net419 vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__mux2_1
X_13391_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] _05705_ vssd1 vssd1
+ vccd1 vccd1 _03852_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08615__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13050__S net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15130_ net1370 vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__inv_2
X_12342_ net2821 net260 net429 vssd1 vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15061_ net1274 vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__inv_2
X_12273_ net2413 net266 net436 vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08918__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14012_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[89\] _04241_ _04244_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[97\]
+ _04293_ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__a221o_1
X_11224_ net523 _07124_ _07563_ vssd1 vssd1 vccd1 vccd1 _07564_ sky130_fd_sc_hd__o21a_1
XFILLER_0_120_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12902__B net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09591__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11155_ _07211_ _07214_ net519 vssd1 vssd1 vccd1 vccd1 _07495_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_147_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10106_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[6\] net743 net732 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06446_ sky130_fd_sc_hd__a22o_1
X_11086_ _05805_ net513 vssd1 vssd1 vccd1 vccd1 _07426_ sky130_fd_sc_hd__nor2_1
X_15963_ net1367 vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_125_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17702_ clknet_leaf_134_wb_clk_i _03386_ _01643_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[23\]
+ sky130_fd_sc_hd__dfrtp_4
X_10037_ net1143 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[0\] net981 vssd1
+ vssd1 vccd1 vccd1 _06377_ sky130_fd_sc_hd__and3_1
X_14914_ net1350 vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__inv_2
X_15894_ net1408 vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__inv_2
XANTENNA__09894__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17633_ clknet_leaf_0_wb_clk_i _03318_ _01574_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_19_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14845_ net1241 vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_121_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17564_ clknet_leaf_88_wb_clk_i _03251_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_14776_ net1217 vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__inv_2
X_11988_ net2034 net306 net474 vssd1 vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09646__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09004__A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08546__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13727_ _03735_ _04098_ vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__nand2_1
X_16515_ clknet_leaf_1_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[13\]
+ _00498_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10939_ _07185_ _07278_ _07276_ vssd1 vssd1 vccd1 vccd1 _07279_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11453__A2 _04621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17495_ clknet_leaf_15_wb_clk_i _03182_ _01478_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10661__A0 _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16446_ clknet_leaf_52_wb_clk_i _02200_ _00429_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_144_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13658_ net187 _04089_ _04090_ net728 vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12609_ net2415 net225 net395 vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__mux2_1
XANTENNA__11205__A2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16377_ clknet_leaf_99_wb_clk_i _02131_ _00360_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[100\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13589_ net198 net194 _07811_ _07883_ net644 vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_26_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10437__X _06777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15328_ net1234 vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_134_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_134_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__15676__A net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15259_ net1274 vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__inv_2
XANTENNA__10316__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09674__A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09820_ net376 _05378_ _05416_ _05454_ net560 vssd1 vssd1 vccd1 vccd1 _06160_ sky130_fd_sc_hd__a41o_1
Xfanout407 _03564_ vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__clkbuf_8
Xfanout418 _03562_ vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__buf_4
XFILLER_0_10_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12304__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout429 _07965_ vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__clkbuf_8
X_09751_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[20\] net815 net753 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__a22o_1
XANTENNA__12469__A1 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08702_ net603 net585 _05041_ vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__a21o_1
XFILLER_0_146_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13130__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09682_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[22\] net807 net787 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__a22o_1
XANTENNA__11141__A1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08542__C1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08633_ net1020 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[10\] net898 vssd1
+ vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout268_A _07877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08564_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[19\] net696 _04901_
+ _04902_ _04903_ vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_89_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14091__B1 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08495_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[23\] net686 _04784_ _04822_
+ net705 vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12827__X _03648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08845__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout435_A net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1177_A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08753__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13197__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout602_A net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1344_A net1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09116_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] _04846_ net593 vssd1 vssd1
+ vccd1 vccd1 _05456_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_17_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09287__C net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09047_ net1111 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[12\] net932
+ vssd1 vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1132_X net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold450 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[0\] vssd1 vssd1 vccd1 vccd1
+ net1985 sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[10\] vssd1 vssd1 vccd1 vccd1
+ net1996 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout971_A _04645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold472 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2007 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10707__B2 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold483 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2018 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold494 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2029 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12214__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10523__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10183__A2 _04678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout930 net933 vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__clkbuf_2
Xfanout941 net942 vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__buf_4
X_09949_ net998 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[3\] net955 vssd1
+ vssd1 vccd1 vccd1 _06289_ sky130_fd_sc_hd__and3_1
Xfanout952 net953 vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout963 _04653_ vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout974 _04640_ vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_70_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13121__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout985 _04629_ vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__buf_4
X_12960_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[2\] _05258_ net1039 vssd1
+ vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__mux2_1
Xfanout996 net997 vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1150 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[35\] vssd1 vssd1 vccd1 vccd1
+ net2685 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11911_ net2526 net256 net480 vssd1 vssd1 vccd1 vccd1 _03068_ sky130_fd_sc_hd__mux2_1
Xhold1161 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2696 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16567__D net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1172 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2707 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12880__A1 _05779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12891_ net2197 net871 net358 _03668_ vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__a22o_1
Xhold1183 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[79\] vssd1 vssd1 vccd1 vccd1
+ net2718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1194 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2729 sky130_fd_sc_hd__dlygate4sd3_1
X_14630_ net1293 vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__inv_2
XANTENNA__11354__A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11842_ net2274 net263 net487 vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__mux2_1
XANTENNA__10891__B1 _07230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09628__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14082__B1 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11073__B _06707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14561_ net1411 vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__inv_2
X_11773_ net1766 net265 net498 vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__mux2_1
XANTENNA__12884__S net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10643__A0 _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11641__X _07851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13512_ net187 _03968_ _03969_ net727 vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__a211o_1
X_16300_ clknet_leaf_120_wb_clk_i _02054_ _00283_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_17280_ clknet_leaf_48_wb_clk_i _02967_ _01263_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10724_ _07061_ _07063_ net517 vssd1 vssd1 vccd1 vccd1 _07064_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14492_ net1406 vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__inv_2
X_16231_ clknet_leaf_130_wb_clk_i net2198 _00219_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__dfrtp_1
XANTENNA__13188__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13443_ _03901_ _03903_ vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__and2_1
X_10655_ net533 _06994_ _06993_ _05263_ vssd1 vssd1 vccd1 vccd1 _06995_ sky130_fd_sc_hd__a211o_1
XANTENNA__11199__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08382__B team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16162_ clknet_leaf_131_wb_clk_i _01925_ _00150_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13374_ net1562 net829 _03838_ team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1
+ vccd1 vccd1 _01873_ sky130_fd_sc_hd__a22o_1
Xclkload17 clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload17/Y sky130_fd_sc_hd__inv_6
XANTENNA__09197__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10586_ net503 _06882_ net333 _06925_ vssd1 vssd1 vccd1 vccd1 _06926_ sky130_fd_sc_hd__a31o_1
Xclkload28 clknet_leaf_148_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload28/Y sky130_fd_sc_hd__inv_6
XANTENNA__09261__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09800__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15113_ net1294 vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__inv_2
Xclkload39 clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload39/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_50_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12325_ net2874 net190 net427 vssd1 vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__mux2_1
X_16093_ clknet_leaf_132_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[15\]
+ _00081_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12913__A _04881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17984__1499 vssd1 vssd1 vccd1 vccd1 _17984__1499/HI net1499 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_114_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15044_ net1233 vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_114_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12256_ net2121 net314 net441 vssd1 vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__mux2_1
X_11207_ _06915_ _07369_ _07371_ net335 _07546_ vssd1 vssd1 vccd1 vccd1 _07547_ sky130_fd_sc_hd__o221a_1
XFILLER_0_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12187_ net2493 net320 net450 vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__mux2_1
XANTENNA__10174__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11138_ _06402_ _06403_ _07477_ vssd1 vssd1 vccd1 vccd1 _07478_ sky130_fd_sc_hd__o21a_1
X_16995_ clknet_leaf_26_wb_clk_i _02682_ _00978_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09316__A1 net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11963__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13112__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11069_ _07408_ _07377_ vssd1 vssd1 vccd1 vccd1 _07409_ sky130_fd_sc_hd__nand2b_1
X_15946_ net1363 vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__inv_2
XANTENNA__09867__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15877_ net1356 vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17616_ clknet_leaf_2_wb_clk_i _03301_ _01557_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_59_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14828_ net1258 vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__inv_2
XANTENNA__13182__C net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14073__B1 _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09619__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17547_ clknet_leaf_5_wb_clk_i _03234_ _01530_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_14759_ net1311 vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08280_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[1\] net1872 net1043 vssd1 vssd1
+ vccd1 vccd1 _03407_ sky130_fd_sc_hd__mux2_1
XANTENNA__09669__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17478_ clknet_leaf_73_wb_clk_i _03165_ _01461_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12807__B _07308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13179__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16429_ clknet_leaf_135_wb_clk_i _02183_ _00412_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08292__B net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12926__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12823__A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08358__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10343__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout204 _07855_ vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__buf_2
XANTENNA__12034__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout215 net217 vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10165__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout226 net228 vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__clkbuf_2
X_09803_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[14\] net802 net778 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[14\]
+ _06136_ vssd1 vssd1 vccd1 vccd1 _06143_ sky130_fd_sc_hd__a221o_1
Xfanout237 net238 vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__clkbuf_2
Xfanout248 _07842_ vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__buf_1
Xfanout259 net260 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__clkbuf_2
X_07995_ team_01_WB.instance_to_wrap.cpu.f0.num\[30\] vssd1 vssd1 vccd1 vccd1 _04493_
+ sky130_fd_sc_hd__inv_2
XANTENNA__13639__B1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout385_A _03570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11873__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_105_Left_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09734_ net995 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[20\] net957 vssd1
+ vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_31_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09858__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09665_ net1136 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[22\] net984
+ vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout552_A _05151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09570__C net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1294_A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08616_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[11\] net684 net670 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09596_ net996 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[24\] net976 vssd1
+ vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__and3_1
XANTENNA__14064__B1 _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08547_ net999 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[19\] net901 vssd1
+ vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout340_X net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout817_A net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout438_X net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08478_ net1001 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[23\] net914
+ vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_46_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09491__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_114_Left_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12209__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout605_X net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10518__A net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10440_ _05737_ _05759_ vssd1 vssd1 vccd1 vccd1 _06780_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08770__X _05110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09243__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08597__A2 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10371_ net377 _06709_ _05566_ vssd1 vssd1 vccd1 vccd1 _06711_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_131_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12110_ net2983 net255 net456 vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__mux2_1
X_13090_ _03713_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[4\] net853 vssd1 vssd1
+ vccd1 vccd1 _02035_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout974_X net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12041_ net2451 net261 net463 vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__mux2_1
XANTENNA__11349__A team_01_WB.instance_to_wrap.cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold280 team_01_WB.instance_to_wrap.a1.ADR_I\[21\] vssd1 vssd1 vccd1 vccd1 net1815
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 team_01_WB.instance_to_wrap.cpu.f0.write_data\[20\] vssd1 vssd1 vccd1 vccd1
+ net1826 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17225__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_123_Left_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11783__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout760 net762 vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout771 _04672_ vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11636__X _07847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15800_ net1218 vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__inv_2
Xfanout782 net784 vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__clkbuf_8
X_16780_ clknet_leaf_16_wb_clk_i _02467_ _00763_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13992_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[80\] _04245_ _04266_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__a22o_1
Xfanout793 _04652_ vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15731_ net1392 vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__inv_2
X_12943_ _05373_ _07757_ _03694_ vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__o21ai_2
XANTENNA__08377__B _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15662_ net1292 vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__inv_2
X_12874_ _05833_ _07752_ net361 vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_68_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17401_ clknet_leaf_103_wb_clk_i _03088_ _01384_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14613_ net1308 vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__inv_2
X_11825_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\] team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\]
+ vssd1 vssd1 vccd1 vccd1 _07946_ sky130_fd_sc_hd__and2b_2
X_15593_ net1295 vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14544_ net1352 vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__inv_2
X_17332_ clknet_leaf_66_wb_clk_i _03019_ _01315_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11756_ net2135 net288 net502 vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09482__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08824__C net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10707_ _05805_ net330 _07044_ net368 _07046_ vssd1 vssd1 vccd1 vccd1 _07047_ sky130_fd_sc_hd__o221a_1
XFILLER_0_153_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14475_ net1418 vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__inv_2
X_17263_ clknet_leaf_33_wb_clk_i _02950_ _01246_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12119__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11687_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] _07808_ vssd1 vssd1
+ vccd1 vccd1 _07887_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17933__1450 vssd1 vssd1 vccd1 vccd1 _17933__1450/HI net1450 sky130_fd_sc_hd__conb_1
XFILLER_0_126_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13426_ _03885_ _03886_ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__or2_1
X_16214_ clknet_leaf_124_wb_clk_i _01974_ _00202_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10638_ _06929_ _06969_ vssd1 vssd1 vccd1 vccd1 _06978_ sky130_fd_sc_hd__or2_1
XANTENNA__08037__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17194_ clknet_leaf_30_wb_clk_i _02881_ _01177_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09234__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload106 clknet_leaf_99_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload106/Y sky130_fd_sc_hd__inv_8
Xclkload117 clknet_leaf_72_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload117/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload128 clknet_leaf_77_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload128/Y sky130_fd_sc_hd__clkinv_8
X_16145_ clknet_leaf_130_wb_clk_i net2486 _00133_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08588__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload139 clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload139/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_144_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10862__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13357_ _04483_ _07684_ vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__nand2_1
X_10569_ _06907_ _06908_ net536 vssd1 vssd1 vccd1 vccd1 _06909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10395__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12308_ net2200 net231 net433 vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__mux2_1
X_16076_ clknet_leaf_153_wb_clk_i _01869_ _00064_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[31\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_122_885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13288_ team_01_WB.instance_to_wrap.cpu.f0.i\[24\] _03746_ _03774_ vssd1 vssd1 vccd1
+ vccd1 _03775_ sky130_fd_sc_hd__o21a_1
X_15027_ net1394 vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_53_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12239_ net2425 net235 net439 vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__mux2_1
XANTENNA__10147__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09952__A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12789__S net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11693__S net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08760__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16978_ clknet_leaf_110_wb_clk_i _02665_ _00961_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput4 DAT_I[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
X_15929_ net1408 vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09450_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[29\] net651 net649 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__a22o_1
XANTENNA__14046__B1 _04230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08401_ _04733_ _04739_ _04740_ vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__and3b_1
XFILLER_0_59_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09381_ net1115 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[26\] net909
+ _04797_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[26\] vssd1 vssd1 vccd1
+ vccd1 _05721_ sky130_fd_sc_hd__a32o_1
XFILLER_0_143_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10870__A3 _06707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12818__A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11281__X _07621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08332_ net991 net945 vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__and2_4
XANTENNA__10706__C_N net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08263_ net2304 net2224 net1052 vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12029__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10338__A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_92_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08194_ net2771 net2756 net1047 vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11868__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1042_A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12780__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13309__C1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09565__C net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11169__A _07269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10138__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11335__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12699__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_X net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07978_ team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1 _04476_
+ sky130_fd_sc_hd__inv_2
XANTENNA__08478__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09717_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[21\] net802 net800 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout934_A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08503__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09648_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[23\] net745 net738 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_48_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10310__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17983__1498 vssd1 vssd1 vccd1 vccd1 _17983__1498/HI net1498 sky130_fd_sc_hd__conb_1
XANTENNA__13831__B net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout722_X net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09579_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[25\] net820 net777 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11632__A net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11610_ _07821_ _07825_ vssd1 vssd1 vccd1 vccd1 _07826_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_26_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ net2660 net223 net395 vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09102__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08644__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11541_ net1662 net1174 net590 net1169 vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10248__A net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14260_ net1205 vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__inv_2
X_11472_ net366 _07763_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[27\] net874
+ vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_151_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11778__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13211_ net28 net836 net629 net1813 vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__o22a_1
X_10423_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[27\] net759 net752 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06763_ sky130_fd_sc_hd__a22o_1
X_14191_ _04458_ _04459_ vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12771__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13142_ net1637 net845 net633 team_01_WB.instance_to_wrap.a1.ADR_I\[1\] vssd1 vssd1
+ vccd1 vccd1 _01999_ sky130_fd_sc_hd__a22o_1
X_10354_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[17\] net760 _06680_
+ _06684_ _06690_ vssd1 vssd1 vccd1 vccd1 _06694_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_111_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input63_A wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_111_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09475__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17950_ net1465 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
XFILLER_0_20_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13073_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[13\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[21\]
+ net860 vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__mux2_1
X_10285_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[19\] net791 net749 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _06625_ sky130_fd_sc_hd__a22o_1
XANTENNA__10414__C net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16901_ clknet_leaf_46_wb_clk_i _02588_ _00884_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12024_ net1787 net291 net470 vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__mux2_1
X_17881_ clknet_leaf_139_wb_clk_i _03556_ _01821_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_16832_ clknet_leaf_46_wb_clk_i _02519_ _00815_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_137_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12402__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout590 _07785_ vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__buf_2
XANTENNA__08819__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16763_ clknet_leaf_70_wb_clk_i _02450_ _00746_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_109_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12826__A1 _07489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13975_ _04217_ _04219_ _04227_ vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__and3_4
X_15714_ net1319 vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__inv_2
X_12926_ net2239 net871 net358 _03693_ vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__a22o_1
X_16694_ clknet_leaf_29_wb_clk_i _02381_ _00677_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15645_ net1315 vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__inv_2
X_12857_ net1954 net301 net382 vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11808_ net2193 net229 net493 vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__mux2_1
X_12788_ net1729 net640 net608 _03620_ vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__a22o_1
X_15576_ net1216 vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09012__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11262__B1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08554__C net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17315_ clknet_leaf_25_wb_clk_i _03002_ _01298_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11739_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\]
+ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] vssd1 vssd1 vccd1 vccd1 _07929_
+ sky130_fd_sc_hd__a21oi_1
X_14527_ net1404 vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17246_ clknet_leaf_85_wb_clk_i _02933_ _01229_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09947__A net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08851__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14458_ net1305 vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_12_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13554__A2 _07621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13469__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09758__B2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13409_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] _05220_ vssd1 vssd1 vccd1
+ vccd1 _03870_ sky130_fd_sc_hd__and2_1
X_17177_ clknet_leaf_72_wb_clk_i _02864_ _01160_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14389_ net1186 vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12762__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16128_ clknet_leaf_126_wb_clk_i _00019_ _00116_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_08950_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[6\] net660 _05272_ _05273_
+ _05289_ vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__a2111o_1
X_16059_ clknet_leaf_154_wb_clk_i _01852_ _00047_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10324__C net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08881_ net602 _05220_ vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_135_Right_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17672__Q team_01_WB.instance_to_wrap.cpu.DM0.readdata\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12312__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12817__B2 _03640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09502_ net1150 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[29\] net977
+ vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__and3_1
XFILLER_0_154_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10828__B1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08448__D net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08497__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[23\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1032 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09433_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[28\] net692 net684 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[28\]
+ _05772_ vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout250_A _07904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09364_ _05691_ _05692_ _05703_ net703 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__o32a_2
XTAP_TAPCELL_ROW_43_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11171__B net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08315_ net1131 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[30\] net963
+ vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_20 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12982__S net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09295_ net1083 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[22\] net925
+ vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_31 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout515_A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1257_A net1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_42 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09857__A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_53 _03654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08246_ net2685 net2587 net1055 vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__mux2_1
XANTENNA_64 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_958 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08177_ net3020 net2956 net1047 vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10359__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12753__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09295__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout884_A net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput160 net160 vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_2
Xoutput171 net171 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__clkbuf_4
Xoutput182 net182 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__clkbuf_4
XANTENNA__09592__A net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10070_ _06406_ _06408_ _06254_ _06285_ vssd1 vssd1 vccd1 vccd1 _06410_ sky130_fd_sc_hd__o211ai_4
XANTENNA_fanout672_X net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13826__B net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11186__X _07526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08724__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09382__C1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12222__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10531__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08639__C net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11346__B team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08001__A net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13744__B1_N net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout937_X net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13760_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[8\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[11\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__and4bb_1
X_10972_ _05301_ net372 vssd1 vssd1 vccd1 vccd1 _07312_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_67_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09685__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13481__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12711_ net2891 net301 net384 vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__mux2_1
X_13691_ team_01_WB.instance_to_wrap.cpu.c0.count\[11\] team_01_WB.instance_to_wrap.cpu.c0.count\[8\]
+ team_01_WB.instance_to_wrap.cpu.c0.count\[7\] team_01_WB.instance_to_wrap.cpu.c0.count\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__or4bb_1
XTAP_TAPCELL_ROW_104_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12642_ net2330 net226 net391 vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__mux2_1
X_15430_ net1380 vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__inv_2
XANTENNA__09437__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15361_ net1279 vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__inv_2
X_12573_ net2275 net257 net401 vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17100_ clknet_leaf_20_wb_clk_i _02787_ _01083_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11795__A1 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11524_ net1705 net1171 net588 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] vssd1
+ vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__a22o_1
X_14312_ net1325 vssd1 vssd1 vccd1 vccd1 _00106_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15292_ net1247 vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14243_ net1236 vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__inv_2
X_17031_ clknet_leaf_107_wb_clk_i _02718_ _01014_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13536__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11455_ net1175 team_01_WB.instance_to_wrap.cpu.DM0.state\[2\] vssd1 vssd1 vccd1
+ vccd1 team_01_WB.instance_to_wrap.cpu.DM0.next_enable sky130_fd_sc_hd__and2_1
XFILLER_0_22_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12744__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10406_ net505 _06638_ _06675_ vssd1 vssd1 vccd1 vccd1 _06746_ sky130_fd_sc_hd__o21bai_1
X_14174_ net2006 _04447_ net1183 vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11386_ team_01_WB.instance_to_wrap.cpu.f0.i\[28\] net1068 _07668_ _07714_ vssd1
+ vssd1 vccd1 vccd1 _07715_ sky130_fd_sc_hd__nand4_2
XFILLER_0_68_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13125_ net84 net843 net631 net1722 vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__a22o_1
X_10337_ _06675_ _06676_ vssd1 vssd1 vccd1 vccd1 _06677_ sky130_fd_sc_hd__nand2_1
X_17933_ net1450 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
X_13056_ net2846 net2765 net853 vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__mux2_1
X_10268_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[19\] net804 _06605_
+ _06606_ _06607_ vssd1 vssd1 vccd1 vccd1 _06608_ sky130_fd_sc_hd__a2111o_1
X_12007_ net3160 net265 net467 vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__mux2_1
Xfanout1330 net1332 vssd1 vssd1 vccd1 vccd1 net1330 sky130_fd_sc_hd__buf_4
XANTENNA__09912__A1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1341 net1343 vssd1 vssd1 vccd1 vccd1 net1341 sky130_fd_sc_hd__buf_4
XANTENNA__10441__A net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17864_ clknet_leaf_125_wb_clk_i _03539_ _01804_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12132__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1352 net1355 vssd1 vssd1 vccd1 vccd1 net1352 sky130_fd_sc_hd__buf_4
XFILLER_0_84_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10199_ net1142 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[8\] net958 vssd1
+ vssd1 vccd1 vccd1 _06539_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_159_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_159_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout1363 net1365 vssd1 vssd1 vccd1 vccd1 net1363 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_128_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1374 net1377 vssd1 vssd1 vccd1 vccd1 net1374 sky130_fd_sc_hd__buf_4
XFILLER_0_17_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1385 net1387 vssd1 vssd1 vccd1 vccd1 net1385 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_128_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16815_ clknet_leaf_35_wb_clk_i _02502_ _00798_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1396 net1397 vssd1 vssd1 vccd1 vccd1 net1396 sky130_fd_sc_hd__clkbuf_4
X_17795_ clknet_leaf_94_wb_clk_i _03471_ _01735_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[65\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14848__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11971__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16746_ clknet_leaf_10_wb_clk_i _02433_ _00729_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09676__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13958_ _04238_ _04248_ vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__nor2_4
XANTENNA__09441__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09140__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12909_ net1641 net869 net356 _03681_ vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__a22o_1
X_16677_ clknet_leaf_52_wb_clk_i _02364_ _00660_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13889_ net1426 _04146_ _04195_ vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__nor3_1
XFILLER_0_146_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15628_ net1259 vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09428__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13224__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_118_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15559_ net1389 vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__inv_2
X_08100_ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[3\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[2\]
+ _04569_ _04570_ vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__or4_1
XFILLER_0_71_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09080_ net1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[13\] net905
+ vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08581__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08031_ net1592 net568 net347 team_01_WB.instance_to_wrap.cpu.f0.i\[24\] vssd1 vssd1
+ vccd1 vccd1 _03560_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16571__Q team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput40 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_1
X_17229_ clknet_leaf_67_wb_clk_i _02916_ _01212_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12307__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12735__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput51 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
Xinput62 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_1
Xhold802 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[103\] vssd1 vssd1 vccd1 vccd1
+ net2337 sky130_fd_sc_hd__dlygate4sd3_1
Xinput73 wbs_stb_i vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11538__B2 net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08453__B_N net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold813 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold824 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[74\] vssd1 vssd1 vccd1 vccd1
+ net2359 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09600__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold835 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[49\] vssd1 vssd1 vccd1 vccd1
+ net2381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2392 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08954__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09982_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[2\] net793 net778 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06322_ sky130_fd_sc_hd__a22o_1
Xhold868 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[105\] vssd1 vssd1 vccd1 vccd1
+ net2403 sky130_fd_sc_hd__dlygate4sd3_1
X_17982__1497 vssd1 vssd1 vccd1 vccd1 _17982__1497/HI net1497 sky130_fd_sc_hd__conb_1
Xhold879 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2414 sky130_fd_sc_hd__dlygate4sd3_1
X_08933_ net1111 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[6\] net912 vssd1
+ vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout298_A _07921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13160__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08864_ net1018 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[3\] net936 vssd1
+ vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__and3_1
Xhold1502 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net3037 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12042__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1513 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3048 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1005_A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1524 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net3059 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1535 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net3070 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1546 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net3081 sky130_fd_sc_hd__dlygate4sd3_1
X_08795_ net1009 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[0\] net914 vssd1
+ vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__and3_1
Xhold1557 team_01_WB.instance_to_wrap.cpu.f0.num\[31\] vssd1 vssd1 vccd1 vccd1 net3092
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14758__A net1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1568 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net3103 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11881__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout465_A _07954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1579 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net3114 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_28_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14110__X _04396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08756__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_2_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13381__B _05803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11474__B1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout632_A _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10816__A3 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08475__B net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09416_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[27\] net701 _05749_ _05755_
+ vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__o22a_1
XFILLER_0_137_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09347_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[25\] _04776_ net685 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout420_X net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13620__D1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout518_X net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09278_ net597 _05615_ _05617_ vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__o21ai_4
XANTENNA__13518__A2 _07566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08229_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[52\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[44\]
+ net1050 vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__mux2_1
XANTENNA__12217__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1427_X net1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11529__B2 net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11240_ _06750_ _06817_ _06822_ net343 vssd1 vssd1 vccd1 vccd1 _07580_ sky130_fd_sc_hd__a31o_1
XFILLER_0_31_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout887_X net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10960__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11171_ _05416_ net330 vssd1 vssd1 vccd1 vccd1 _07511_ sky130_fd_sc_hd__nor2_1
X_10122_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[6\] net778 net747 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06462_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13151__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14930_ net1292 vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__inv_2
X_10053_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[0\] net824 net794 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06393_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11701__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10504__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input26_A DAT_I[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09370__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14861_ net1261 vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__inv_2
XANTENNA__12887__S net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16600_ clknet_leaf_49_wb_clk_i _02287_ _00583_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13812_ net2917 net833 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[5\]
+ sky130_fd_sc_hd__and2_1
X_17580_ clknet_leaf_95_wb_clk_i _03267_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__dfxtp_1
X_14792_ net1375 vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_123_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16531_ clknet_leaf_159_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[29\]
+ _00514_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_123_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13743_ _04136_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__inv_2
X_10955_ _05043_ _06438_ vssd1 vssd1 vccd1 vccd1 _07295_ sky130_fd_sc_hd__nor2_1
XANTENNA__11092__A net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16462_ clknet_leaf_113_wb_clk_i _02216_ _00445_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13674_ net1584 net567 net345 net1068 vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__a22o_1
X_10886_ net327 _07219_ _07221_ _07225_ vssd1 vssd1 vccd1 vccd1 _07226_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_14_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15413_ net1285 vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12625_ net2044 net215 net392 vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__mux2_1
X_16393_ clknet_leaf_97_wb_clk_i _02147_ _00376_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[116\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_81_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09497__A _04706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12965__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12556_ net2998 net190 net399 vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15344_ net1279 vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14167__C1 net1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11507_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[9\] _07756_ vssd1 vssd1 vccd1
+ vccd1 _07781_ sky130_fd_sc_hd__and2_1
XANTENNA__08832__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15275_ net1395 vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__inv_2
X_12487_ net2007 net313 net413 vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__mux2_1
XANTENNA__12127__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold109 net97 vssd1 vssd1 vccd1 vccd1 net1644 sky130_fd_sc_hd__dlygate4sd3_1
X_17014_ clknet_leaf_12_wb_clk_i _02701_ _00997_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11438_ _07736_ _07743_ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__nor2_1
X_14226_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[6\] vssd1 vssd1 vccd1
+ vccd1 _02261_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_145_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13857__A_N net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11966__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14157_ _04195_ _04438_ net1421 vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__a21oi_1
X_11369_ _07670_ _07697_ vssd1 vssd1 vccd1 vccd1 _07698_ sky130_fd_sc_hd__nand2_1
X_13108_ team_01_WB.EN_VAL_REG net72 _03730_ vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__mux2_1
X_14088_ _04348_ _04375_ _04356_ net1183 vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__o211a_1
XANTENNA__09663__C net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13142__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17916_ net1523 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
X_13039_ net2836 net2757 net856 vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1160 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[18\] vssd1 vssd1 vccd1 vccd1
+ net1160 sky130_fd_sc_hd__clkbuf_2
Xfanout1171 net1172 vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__buf_2
XANTENNA__09361__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17847_ clknet_leaf_98_wb_clk_i _03523_ _01787_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[117\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout1193 net1201 vssd1 vssd1 vccd1 vccd1 net1193 sky130_fd_sc_hd__buf_4
XFILLER_0_156_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08580_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[15\] net680 net647 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__a22o_1
X_17778_ clknet_leaf_123_wb_clk_i net2617 _01718_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09113__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16566__Q team_01_WB.instance_to_wrap.cpu.DM0.dhit vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16729_ clknet_leaf_102_wb_clk_i _02416_ _00712_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09201_ net1087 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[17\] net929
+ vssd1 vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_56_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09132_ net1024 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[14\] net927 vssd1
+ vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08742__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09063_ net1111 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[12\] net928
+ vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__and3_1
X_17895__1517 vssd1 vssd1 vccd1 vccd1 net1517 _17895__1517/LO sky130_fd_sc_hd__conb_1
XFILLER_0_72_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12037__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10346__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout213_A _07838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08014_ team_01_WB.instance_to_wrap.cpu.RU0.state\[0\] vssd1 vssd1 vccd1 vccd1 _04510_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_114_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold610 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2145 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold621 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2156 sky130_fd_sc_hd__dlygate4sd3_1
Xhold632 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2167 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11876__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold643 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 net2178
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11729__X _07921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold654 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2189 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold665 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold676 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold687 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[50\] vssd1 vssd1 vccd1 vccd1
+ net2222 sky130_fd_sc_hd__dlygate4sd3_1
Xhold698 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2233 sky130_fd_sc_hd__dlygate4sd3_1
X_09965_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[3\] net823 _06287_ _06290_
+ _06296_ vssd1 vssd1 vccd1 vccd1 _06305_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08103__X _04574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09573__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08916_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[2\] net672 _05226_ _05228_
+ _05233_ vssd1 vssd1 vccd1 vccd1 _05256_ sky130_fd_sc_hd__a2111o_1
X_09896_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[5\] net809 _06223_ _06224_
+ _06231_ vssd1 vssd1 vccd1 vccd1 _06236_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout1008_X net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1310 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2845 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_86_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1321 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[35\] vssd1 vssd1 vccd1 vccd1
+ net2856 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09352__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1332 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2867 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout370_X net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1343 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[86\] vssd1 vssd1 vccd1 vccd1
+ net2878 sky130_fd_sc_hd__dlygate4sd3_1
X_08847_ _05178_ _05182_ _05186_ _05155_ vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__o31a_4
XANTENNA__17860__Q team_01_WB.instance_to_wrap.cpu.RU0.InstrRead vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold1354 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2889 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout847_A net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout468_X net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13392__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1365 team_01_WB.instance_to_wrap.cpu.f0.num\[18\] vssd1 vssd1 vccd1 vccd1 net2900
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1376 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2911 sky130_fd_sc_hd__dlygate4sd3_1
X_08778_ net1010 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[0\] net917 vssd1
+ vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__and3_1
Xhold1387 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2922 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12500__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1398 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2933 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09104__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13987__A2 _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_3_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10740_ _06982_ _06999_ net533 vssd1 vssd1 vccd1 vccd1 _07080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout802_X net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10671_ _07010_ vssd1 vssd1 vccd1 vccd1 _07011_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12410_ net3046 net287 net421 vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__mux2_1
XANTENNA__11640__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13390_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] _05705_ vssd1 vssd1
+ vccd1 vccd1 _03851_ sky130_fd_sc_hd__or2_1
XANTENNA__09812__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10958__C1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08652__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14149__C1 _04152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12341_ net2939 net231 net429 vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15060_ net1379 vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_79_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12272_ net2740 net235 net435 vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11786__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14011_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[41\] _04246_ _04261_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[113\]
+ _04292_ vssd1 vssd1 vccd1 vccd1 _04302_ sky130_fd_sc_hd__a221o_1
XANTENNA__08918__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11223_ _06890_ _06906_ _06909_ _05263_ net338 vssd1 vssd1 vccd1 vccd1 _07563_ sky130_fd_sc_hd__o221a_1
XFILLER_0_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09040__A1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09591__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11154_ net344 _07492_ _07493_ vssd1 vssd1 vccd1 vccd1 _07494_ sky130_fd_sc_hd__or3_1
XFILLER_0_101_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10105_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[6\] net823 net796 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[6\]
+ _06443_ vssd1 vssd1 vccd1 vccd1 _06445_ sky130_fd_sc_hd__a221o_1
XFILLER_0_105_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11085_ _05759_ net504 _07347_ _07423_ _07424_ vssd1 vssd1 vccd1 vccd1 _07425_ sky130_fd_sc_hd__o221a_1
X_15962_ net1363 vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__inv_2
XANTENNA__13675__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17701_ clknet_leaf_134_wb_clk_i _03385_ _01642_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10422__C net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10036_ net1142 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[0\] net948 vssd1
+ vssd1 vccd1 vccd1 _06376_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_125_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14913_ net1279 vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_125_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11686__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15893_ net1415 vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17632_ clknet_leaf_3_wb_clk_i _03317_ _01573_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12410__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14844_ net1246 vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08827__C net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17563_ clknet_leaf_89_wb_clk_i _03250_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13978__A2 _04244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08839__D1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14775_ net1217 vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__inv_2
X_11987_ net2426 net309 net472 vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16514_ clknet_leaf_2_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[12\]
+ _00497_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13726_ net1175 team_01_WB.instance_to_wrap.cpu.f0.state\[7\] _04575_ vssd1 vssd1
+ vccd1 vccd1 _00018_ sky130_fd_sc_hd__a21o_1
XANTENNA__10110__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10938_ net522 _07277_ vssd1 vssd1 vccd1 vccd1 _07278_ sky130_fd_sc_hd__nand2_1
X_17494_ clknet_leaf_12_wb_clk_i _03181_ _01477_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_17981__1496 vssd1 vssd1 vccd1 vccd1 _17981__1496/HI net1496 sky130_fd_sc_hd__conb_1
XFILLER_0_14_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10661__A1 _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16445_ clknet_leaf_45_wb_clk_i _02199_ _00428_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10869_ _06715_ _06740_ _07112_ vssd1 vssd1 vccd1 vccd1 _07209_ sky130_fd_sc_hd__nand3_1
X_13657_ net199 net195 _07934_ net645 vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__o211a_1
XFILLER_0_143_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12608_ net2552 net287 net398 vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__mux2_1
XANTENNA__08606__A1 net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16376_ clknet_leaf_97_wb_clk_i _02130_ _00359_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[99\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09803__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13588_ _03901_ _04032_ vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_30_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08562__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15327_ net1311 vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__inv_2
X_12539_ net1893 net232 net404 vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09955__A net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15258_ net1371 vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13363__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08909__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14209_ net2931 vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15189_ net1282 vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout408 _03564_ vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09582__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout419 net422 vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_103_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_103_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13115__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09750_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[20\] net807 net795 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _06090_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_33_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08701_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] net596 net601 vssd1 vssd1
+ vccd1 vccd1 _05041_ sky130_fd_sc_hd__a21oi_2
XANTENNA__09334__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09681_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[22\] net821 net768 _06011_
+ _06014_ vssd1 vssd1 vccd1 vccd1 _06021_ sky130_fd_sc_hd__a2111o_1
XANTENNA__17680__Q team_01_WB.instance_to_wrap.cpu.f0.i\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08632_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[10\] net912
+ vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__and3_1
XANTENNA__12320__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08737__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08563_ net1077 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[19\] net883
+ vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_81_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08494_ _04830_ _04831_ _04832_ _04833_ vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__or4_1
XFILLER_0_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout330_A _06924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout428_A _07965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09568__C net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09115_ _05454_ vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__inv_2
XANTENNA__08472__C net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1337_A net1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09046_ net1111 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[12\] net893
+ vssd1 vssd1 vccd1 vccd1 _05386_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13354__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13387__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold440 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1975 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10804__A _06919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold451 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1986 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10707__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09076__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold462 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1997 sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2008 sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2019 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold495 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[7\] vssd1 vssd1 vccd1 vccd1
+ net2030 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout964_A _04653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout920 net921 vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__clkbuf_4
Xfanout931 net932 vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__clkbuf_4
Xfanout942 _04759_ vssd1 vssd1 vccd1 vccd1 net942 sky130_fd_sc_hd__buf_4
X_09948_ net1156 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[3\] net949 vssd1
+ vssd1 vccd1 vccd1 _06288_ sky130_fd_sc_hd__and3_1
Xfanout953 _04662_ vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout964 _04653_ vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout975 net976 vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__buf_4
Xfanout986 net987 vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09325__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13834__B net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout752_X net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09879_ net341 _06217_ vssd1 vssd1 vccd1 vccd1 _06219_ sky130_fd_sc_hd__nand2b_1
Xfanout997 net998 vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_142_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1140 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[65\] vssd1 vssd1 vccd1 vccd1
+ net2675 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_142_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1151 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2686 sky130_fd_sc_hd__dlygate4sd3_1
X_11910_ net3070 net259 net481 vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__mux2_1
Xhold1162 team_01_WB.instance_to_wrap.cpu.f0.num\[17\] vssd1 vssd1 vccd1 vccd1 net2697
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12230__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1173 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2708 sky130_fd_sc_hd__dlygate4sd3_1
X_12890_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[25\] _03667_ net1039 vssd1
+ vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__mux2_1
XANTENNA__12880__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1184 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2719 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1195 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[94\] vssd1 vssd1 vccd1 vccd1
+ net2730 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08647__C net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10891__A1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11841_ net2203 net266 net487 vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__mux2_1
X_14560_ net1352 vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__inv_2
X_11772_ net2022 net234 net495 vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10643__A1 _06707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13511_ net198 net194 _07834_ net644 vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__o211a_1
X_10723_ _07062_ vssd1 vssd1 vccd1 vccd1 _07063_ sky130_fd_sc_hd__inv_2
X_14491_ net1415 vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16230_ clknet_leaf_135_wb_clk_i _01990_ _00218_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__dfrtp_1
X_10654_ _05898_ net504 net543 vssd1 vssd1 vccd1 vccd1 _06994_ sky130_fd_sc_hd__mux2_1
X_13442_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] _05456_ vssd1 vssd1
+ vccd1 vccd1 _03903_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16161_ clknet_leaf_134_wb_clk_i _01924_ _00149_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13373_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[6\] net829 _03838_ team_01_WB.instance_to_wrap.cpu.f0.i\[4\]
+ vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10585_ _06882_ net331 _06922_ vssd1 vssd1 vccd1 vccd1 _06925_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_36_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload18 clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload18/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload29 clknet_leaf_149_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload29/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_77_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15112_ net1392 vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_77_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10417__C net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12324_ _07790_ _07794_ net574 vssd1 vssd1 vccd1 vccd1 _07965_ sky130_fd_sc_hd__and3_4
X_16092_ clknet_leaf_132_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[14\]
+ _00080_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[14\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_1_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_51_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12913__B net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12255_ net3143 net319 net442 vssd1 vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__mux2_1
X_15043_ net1270 vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_43_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12405__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10159__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10714__A net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11206_ _05455_ _07545_ vssd1 vssd1 vccd1 vccd1 _07546_ sky130_fd_sc_hd__nand2_1
X_12186_ net2259 net306 net450 vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__mux2_1
X_11137_ _06402_ _06403_ net344 vssd1 vssd1 vccd1 vccd1 _07477_ sky130_fd_sc_hd__a21oi_1
X_16994_ clknet_leaf_57_wb_clk_i _02681_ _00977_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13648__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09316__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11068_ _05338_ _06562_ _07259_ net339 _05374_ vssd1 vssd1 vccd1 vccd1 _07408_ sky130_fd_sc_hd__o32a_1
X_15945_ net1403 vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10019_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[1\] net788 net731 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[1\]
+ _06344_ vssd1 vssd1 vccd1 vccd1 _06359_ sky130_fd_sc_hd__a221o_1
XANTENNA__12140__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17894__1516 vssd1 vssd1 vccd1 vccd1 net1516 _17894__1516/LO sky130_fd_sc_hd__conb_1
XANTENNA__10331__B1 _06669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15876_ net1362 vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__inv_2
XANTENNA__09015__A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17615_ clknet_leaf_2_wb_clk_i _03300_ _01556_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08557__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14827_ net1424 vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17546_ clknet_leaf_31_wb_clk_i _03233_ _01529_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_14758_ net1383 vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__inv_2
XANTENNA__08854__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13709_ _04100_ _04124_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[1\]
+ sky130_fd_sc_hd__and2_1
X_17477_ clknet_leaf_51_wb_clk_i _03164_ _01460_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_14689_ net1205 vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16428_ clknet_leaf_140_wb_clk_i _02182_ _00411_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_82_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_15_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16359_ clknet_leaf_91_wb_clk_i net2803 _00342_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[82\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09252__A1 net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10398__A0 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14128__A2 _04245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17675__Q team_01_WB.instance_to_wrap.cpu.DM0.readdata\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12315__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09555__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout205 _07855_ vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__buf_2
Xfanout216 net217 vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__buf_2
X_09802_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[14\] net757 net753 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[14\]
+ _06137_ vssd1 vssd1 vccd1 vccd1 _06142_ sky130_fd_sc_hd__a221o_1
Xfanout227 net228 vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__buf_2
Xfanout238 net240 vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__buf_2
Xfanout249 _07904_ vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__buf_2
XANTENNA__10911__X _07251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07994_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1 vccd1 _04492_
+ sky130_fd_sc_hd__inv_2
XANTENNA__13639__A1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09307__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09733_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[20\] net779 net752 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _06073_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout280_A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11455__A net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12050__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09664_ net1144 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[22\] net973
+ vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__and3_1
XANTENNA__08467__C net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13941__Y _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08615_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[11\] net688 net679 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[11\]
+ _04953_ vssd1 vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09595_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[24\] net822 net798 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_71_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08546_ net999 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[19\] net935 vssd1
+ vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11461__Y _07757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08477_ net1031 net915 vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout333_X net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08483__B net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09298__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire617 _05335_ vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout500_X net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08046__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1242_X net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_149_Right_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10370_ net377 _05566_ _06709_ vssd1 vssd1 vccd1 vccd1 _06710_ sky130_fd_sc_hd__and3_1
XANTENNA__14119__A2 _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13829__B net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08930__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09029_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[9\] net661 _05346_ _05356_
+ _05357_ vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_131_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10421__A_N net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12040_ net1781 net268 net463 vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold270 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[11\] vssd1 vssd1 vccd1 vccd1
+ net1805 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_72_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09546__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold281 team_01_WB.instance_to_wrap.cpu.c0.count\[10\] vssd1 vssd1 vccd1 vccd1 net1816
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1827 sky130_fd_sc_hd__dlygate4sd3_1
X_17980__1495 vssd1 vssd1 vccd1 vccd1 _17980__1495/HI net1495 sky130_fd_sc_hd__conb_1
XFILLER_0_102_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_127_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout750 _04680_ vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__buf_4
Xfanout761 net762 vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__clkbuf_8
Xfanout772 net774 vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__clkbuf_8
Xfanout783 net784 vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__clkbuf_8
X_13991_ _04279_ _04280_ _04281_ _04282_ vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__or4_1
Xfanout794 net797 vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13056__S net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15730_ net1266 vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__inv_2
X_12942_ _03655_ _03703_ _03704_ net873 net3014 vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__a32o_1
XANTENNA__11084__B _06811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15661_ net1268 vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__inv_2
X_12873_ net1849 net872 net359 _03656_ vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__a22o_1
X_17400_ clknet_leaf_49_wb_clk_i _03087_ _01383_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14612_ net1305 vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__inv_2
X_11824_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\] team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\]
+ vssd1 vssd1 vccd1 vccd1 _07945_ sky130_fd_sc_hd__and2_2
X_15592_ net1398 vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17331_ clknet_leaf_23_wb_clk_i _03018_ _01314_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_14543_ net1406 vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__inv_2
X_11755_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] _07940_ net616 vssd1
+ vssd1 vccd1 vccd1 _07941_ sky130_fd_sc_hd__mux2_2
XANTENNA__09482__A1 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10092__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17262_ clknet_leaf_37_wb_clk_i _02949_ _01245_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11077__A_N net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10706_ _05805_ _06919_ net513 vssd1 vssd1 vccd1 vccd1 _07046_ sky130_fd_sc_hd__or3b_1
X_14474_ net1356 vssd1 vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__inv_2
X_11686_ net719 _07188_ net615 _07885_ vssd1 vssd1 vccd1 vccd1 _07886_ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16213_ clknet_leaf_124_wb_clk_i net1690 _00201_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13425_ _04949_ _03884_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] vssd1
+ vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__o21a_1
XFILLER_0_153_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09001__C net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17193_ clknet_leaf_39_wb_clk_i _02880_ _01176_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10637_ _05835_ _06924_ _06976_ net368 vssd1 vssd1 vccd1 vccd1 _06977_ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload107 clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload107/Y sky130_fd_sc_hd__inv_8
XFILLER_0_102_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload118 clknet_leaf_103_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload118/Y sky130_fd_sc_hd__inv_6
XFILLER_0_24_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload129 clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload129/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16144_ clknet_leaf_128_wb_clk_i _01907_ _00132_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10568_ net504 _06811_ net543 vssd1 vssd1 vccd1 vccd1 _06908_ sky130_fd_sc_hd__mux2_1
X_13356_ _07677_ _03827_ vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12307_ net2309 net264 net433 vssd1 vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__mux2_1
X_16075_ clknet_leaf_156_wb_clk_i _01868_ _00063_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__12135__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13287_ team_01_WB.instance_to_wrap.cpu.f0.i\[24\] _03746_ _04518_ vssd1 vssd1 vccd1
+ vccd1 _03774_ sky130_fd_sc_hd__a21oi_1
X_10499_ net1131 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[31\] net948
+ vssd1 vssd1 vccd1 vccd1 _06839_ sky130_fd_sc_hd__and3b_1
XFILLER_0_122_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15026_ net1290 vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__inv_2
X_12238_ net3034 net237 net439 vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11974__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10552__A0 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12169_ net2986 _07866_ net447 vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09671__C _04662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16977_ clknet_leaf_113_wb_clk_i _02664_ _00960_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput5 DAT_I[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
X_15928_ net1401 vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__inv_2
XANTENNA__10304__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15859_ net1356 vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__inv_2
X_08400_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] _04727_ vssd1 vssd1 vccd1
+ vccd1 _04740_ sky130_fd_sc_hd__nand2_1
X_09380_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[26\] net653 net651 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[26\]
+ _05719_ vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__a221o_1
XANTENNA__08584__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12818__B _07449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16574__Q team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08331_ net1159 net1162 net1165 net1166 vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__nor4_1
XANTENNA_clkbuf_3_7_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17529_ clknet_leaf_71_wb_clk_i _03216_ _01512_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10083__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08262_ net2974 net2847 net1055 vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09225__A1 net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08193_ net2876 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[80\] net1046 vssd1 vssd1
+ vccd1 vccd1 _03494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09776__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08750__C net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12780__A1 _07541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12045__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1035_A team_01_WB.instance_to_wrap.cpu.RU0.InstrRead vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11169__B _07290_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11884__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12532__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout495_A net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08759__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11456__Y _07752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout283_X net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07977_ team_01_WB.instance_to_wrap.cpu.f0.i\[19\] vssd1 vssd1 vccd1 vccd1 _04475_
+ sky130_fd_sc_hd__inv_2
XANTENNA_fanout662_A _04808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13952__X _04244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09716_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[21\] net822 net775 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout450_X net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09647_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[23\] net804 net755 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__a22o_1
XANTENNA__14037__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout927_A net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09578_ _05915_ _05916_ _05917_ vssd1 vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_26_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11191__Y _07531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11632__B _07579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08529_ net1077 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[18\] net901
+ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout715_X net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11540_ net1993 net1174 net590 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1
+ vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13548__B1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11471_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[27\] net579 vssd1 vssd1 vccd1
+ vccd1 _07763_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_154_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13210_ net29 net838 net630 net2917 vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__a22o_1
X_10422_ net1133 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[27\] net964
+ vssd1 vssd1 vccd1 vccd1 _06762_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14190_ net2025 _04457_ net1183 vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17893__1515 vssd1 vssd1 vccd1 vccd1 net1515 _17893__1515/LO sky130_fd_sc_hd__conb_1
XANTENNA__12771__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10353_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[17\] net808 _06679_
+ _06685_ _06689_ vssd1 vssd1 vccd1 vccd1 _06693_ sky130_fd_sc_hd__a2111o_1
X_13141_ net1644 net846 net634 team_01_WB.instance_to_wrap.a1.ADR_I\[2\] vssd1 vssd1
+ vccd1 vccd1 _02000_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_111_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13072_ net2620 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[22\] net853 vssd1 vssd1
+ vccd1 vccd1 _02053_ sky130_fd_sc_hd__mux2_1
XANTENNA__09519__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input56_A wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10284_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[19\] net779 net768 vssd1
+ vssd1 vccd1 vccd1 _06624_ sky130_fd_sc_hd__a21o_1
X_16900_ clknet_leaf_84_wb_clk_i _02587_ _00883_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_12023_ net2204 net315 net469 vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__mux2_1
XANTENNA__11794__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17880_ clknet_leaf_139_wb_clk_i _03555_ _01820_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10534__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16831_ clknet_leaf_41_wb_clk_i _02518_ _00814_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout580 _07752_ vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__clkbuf_2
X_16762_ clknet_leaf_79_wb_clk_i _02449_ _00745_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_109_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13974_ _04217_ _04227_ _04239_ vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__and3_4
X_15713_ net1281 vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__inv_2
X_12925_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[15\] _03692_ net1039 vssd1
+ vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__mux2_1
X_16693_ clknet_leaf_112_wb_clk_i _02380_ _00676_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_15644_ net1253 vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__inv_2
X_12856_ net2412 net281 net381 vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11807_ net1933 net261 net492 vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15575_ net1249 vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__inv_2
X_12787_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] net1062 net365 _03619_
+ vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17314_ clknet_leaf_77_wb_clk_i _03001_ _01297_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14526_ net1351 vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11738_ net716 _07449_ net613 vssd1 vssd1 vccd1 vccd1 _07928_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11969__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17245_ clknet_leaf_64_wb_clk_i _02932_ _01228_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14457_ net1306 vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11669_ _07871_ _07872_ net611 vssd1 vssd1 vccd1 vccd1 _07873_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13408_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] _05112_ vssd1 vssd1 vccd1
+ vccd1 _03869_ sky130_fd_sc_hd__and2_1
XFILLER_0_141_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17176_ clknet_leaf_60_wb_clk_i _02863_ _01159_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09666__C net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14388_ net1188 vssd1 vssd1 vccd1 vccd1 _00182_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08570__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16127_ clknet_leaf_127_wb_clk_i _00018_ _00115_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13339_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[16\] _03814_ net827 vssd1 vssd1
+ vccd1 vccd1 _01884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16058_ clknet_leaf_4_wb_clk_i _01851_ _00046_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_51_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15009_ net1279 vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__inv_2
X_08880_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\] net729 _05111_ net1118 vssd1
+ vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__a22o_2
XANTENNA__09930__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10340__C net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09501_ net1150 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[29\] net952
+ vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_142_Left_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08497__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11733__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09432_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[28\] net697 net675 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08745__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09203__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09363_ _05693_ _05696_ _05700_ _05702_ vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_23_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08314_ net1144 net963 vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_43_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09997__A2 _04678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09294_ net1084 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[22\] net910
+ vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__and3_1
XANTENNA_10 _03663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_21 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_32 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11879__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_43 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08245_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[36\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[28\]
+ net1045 vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__mux2_1
XANTENNA_54 _03654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10783__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout410_A _03564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_65 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1152_A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout508_A _06065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08176_ net2403 net2457 net1056 vssd1 vssd1 vccd1 vccd1 _03511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08480__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1038_X net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput150 net150 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
Xoutput161 net161 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout877_A team_01_WB.instance_to_wrap.cpu.DM0.next_enable vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xoutput172 net172 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout498_X net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput183 net183 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__clkbuf_4
XANTENNA__12503__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1205_X net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09382__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09921__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout665_X net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08776__X _05116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10971_ _06920_ _07141_ _07151_ _06928_ vssd1 vssd1 vccd1 vccd1 _07311_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout832_X net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08488__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12710_ net1961 net280 net384 vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__mux2_1
X_13690_ team_01_WB.instance_to_wrap.cpu.c0.count\[14\] team_01_WB.instance_to_wrap.cpu.c0.count\[13\]
+ team_01_WB.instance_to_wrap.cpu.c0.count\[12\] team_01_WB.instance_to_wrap.cpu.c0.count\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__or4b_1
XFILLER_0_97_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_104_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12641_ net2994 net287 net393 vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_156_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_156_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10047__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11244__A1 _06906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15360_ net1234 vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_156_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09988__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11244__B2 _05263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12572_ net2524 net229 net401 vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11789__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14311_ net1324 vssd1 vssd1 vccd1 vccd1 _00105_ sky130_fd_sc_hd__inv_2
X_11523_ net1629 net1171 net588 team_01_WB.instance_to_wrap.cpu.CU0.bit30 vssd1 vssd1
+ vccd1 vccd1 _03329_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10546__X _06886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15291_ net1254 vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__inv_2
XANTENNA__08660__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17030_ clknet_leaf_90_wb_clk_i _02717_ _01013_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14242_ net1236 vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__inv_2
X_11454_ _07671_ net324 _07751_ vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__and3b_1
XFILLER_0_33_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10706__B _06919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12744__A1 _07566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10405_ _06713_ _06740_ _06712_ vssd1 vssd1 vccd1 vccd1 _06745_ sky130_fd_sc_hd__o21a_1
X_14173_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[8\] _04447_ vssd1 vssd1 vccd1
+ vccd1 _04448_ sky130_fd_sc_hd__and2_1
X_11385_ _04471_ _07713_ vssd1 vssd1 vccd1 vccd1 _07714_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13124_ net1626 net844 net632 team_01_WB.instance_to_wrap.a1.ADR_I\[19\] vssd1 vssd1
+ vccd1 vccd1 _02017_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10336_ _06672_ _06673_ _06674_ vssd1 vssd1 vccd1 vccd1 _06676_ sky130_fd_sc_hd__nand3_1
X_17932_ net1449 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
XANTENNA__12413__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10267_ net990 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[19\] net948 vssd1
+ vssd1 vccd1 vccd1 _06607_ sky130_fd_sc_hd__and3_1
X_13055_ net2769 net2602 net857 vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__mux2_1
XANTENNA__10722__A net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1320 net1321 vssd1 vssd1 vccd1 vccd1 net1320 sky130_fd_sc_hd__buf_4
X_12006_ net2698 net235 net467 vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1331 net1332 vssd1 vssd1 vccd1 vccd1 net1331 sky130_fd_sc_hd__clkbuf_4
X_17863_ clknet_leaf_125_wb_clk_i _03538_ _01803_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10198_ net1139 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[8\] net973 vssd1
+ vssd1 vccd1 vccd1 _06538_ sky130_fd_sc_hd__and3_1
Xfanout1342 net1343 vssd1 vssd1 vccd1 vccd1 net1342 sky130_fd_sc_hd__buf_4
Xfanout1353 net1355 vssd1 vssd1 vccd1 vccd1 net1353 sky130_fd_sc_hd__clkbuf_4
Xfanout1364 net1365 vssd1 vssd1 vccd1 vccd1 net1364 sky130_fd_sc_hd__buf_4
Xfanout1375 net1377 vssd1 vssd1 vccd1 vccd1 net1375 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_128_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16814_ clknet_leaf_27_wb_clk_i _02501_ _00797_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_128_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1386 net1387 vssd1 vssd1 vccd1 vccd1 net1386 sky130_fd_sc_hd__buf_2
X_17794_ clknet_leaf_123_wb_clk_i _03470_ _01734_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[64\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1397 net1398 vssd1 vssd1 vccd1 vccd1 net1397 sky130_fd_sc_hd__buf_4
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16745_ clknet_leaf_39_wb_clk_i _02432_ _00728_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13957_ _04225_ _04248_ vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__nor2_4
XFILLER_0_88_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12908_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[20\] _03680_ net1037 vssd1
+ vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__mux2_1
X_16676_ clknet_leaf_84_wb_clk_i _02363_ _00659_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13888_ _04189_ _04194_ vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__nand2_2
Xclkbuf_leaf_128_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_128_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_33_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15627_ net1424 vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__inv_2
X_12839_ net2015 net246 net380 vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11235__A1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09979__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15558_ net1404 vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__inv_2
XANTENNA__11235__B2 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08862__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11699__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14509_ net1410 vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15489_ net1280 vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__inv_2
X_08030_ team_01_WB.instance_to_wrap.cpu.K0.keyvalid _04523_ _04525_ vssd1 vssd1 vccd1
+ vccd1 _04526_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17228_ clknet_leaf_20_wb_clk_i _02915_ _01211_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput30 DAT_I[6] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
Xinput41 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_1
Xinput52 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12735__A1 _07019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput63 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__clkbuf_1
Xhold803 _02142_ vssd1 vssd1 vccd1 vccd1 net2338 sky130_fd_sc_hd__dlygate4sd3_1
Xinput74 wbs_we_i vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold814 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2349 sky130_fd_sc_hd__dlygate4sd3_1
X_17159_ clknet_leaf_100_wb_clk_i _02846_ _01142_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold825 _03480_ vssd1 vssd1 vccd1 vccd1 net2360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold836 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2371 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold847 _03455_ vssd1 vssd1 vccd1 vccd1 net2382 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09693__A _05657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold858 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2393 sky130_fd_sc_hd__dlygate4sd3_1
X_09981_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[2\] net820 net784 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06321_ sky130_fd_sc_hd__a22o_1
Xhold869 _03519_ vssd1 vssd1 vccd1 vccd1 net2404 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17683__Q team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08932_ net1112 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[6\] net942 vssd1
+ vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__and3_1
XANTENNA__11728__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12323__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09364__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09903__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1503 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[65\] vssd1 vssd1 vccd1 vccd1
+ net3038 sky130_fd_sc_hd__dlygate4sd3_1
X_08863_ net1024 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[3\] net902 vssd1
+ vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_36_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout193_A _07634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1514 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net3049 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1525 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net3060 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_150_Left_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1536 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net3071 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1547 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[8\] vssd1 vssd1 vccd1 vccd1
+ net3082 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_88_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08794_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[0\] net934 vssd1
+ vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__and3_1
Xhold1558 _01931_ vssd1 vssd1 vccd1 vccd1 net3093 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1569 team_01_WB.instance_to_wrap.cpu.c0.count\[6\] vssd1 vssd1 vccd1 vccd1 net3104
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_28_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout360_A net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout458_A _07956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17892__1514 vssd1 vssd1 vccd1 vccd1 net1514 _17892__1514/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_84_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09415_ _05751_ _05752_ _05753_ _05754_ vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_62_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout625_A net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11226__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09346_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[25\] net692 net675 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09277_ net600 _05616_ vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__or2_2
XANTENNA_fanout413_X net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1155_X net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14176__B1 net1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08228_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[53\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[45\]
+ net1053 vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout994_A net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11529__A2 net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08159_ net1672 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[114\] net1052 vssd1 vssd1
+ vccd1 vccd1 _03528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1322_X net1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11170_ _06220_ _07172_ vssd1 vssd1 vccd1 vccd1 _07510_ sky130_fd_sc_hd__nand2_1
XANTENNA__13837__B net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout782_X net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10813__Y _07153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10121_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[6\] net800 _06458_ _06460_
+ vssd1 vssd1 vccd1 vccd1 _06461_ sky130_fd_sc_hd__a211o_1
XFILLER_0_101_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11638__A net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12233__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09355__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10052_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[0\] net730 _06371_ _06372_
+ _06376_ vssd1 vssd1 vccd1 vccd1 _06392_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11162__B1 _07042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11701__A2 _07207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11925__X _07950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14860_ net1257 vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16135__CLK clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13811_ net1813 net833 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[4\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__14100__B1 _04259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14791_ net1389 vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__inv_2
XANTENNA_input19_A DAT_I[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10688__S net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13064__S net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16530_ clknet_leaf_157_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[28\]
+ _00513_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_13742_ net1172 net1032 vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__and2b_1
XANTENNA__10268__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10954_ _07292_ _07293_ vssd1 vssd1 vccd1 vccd1 _07294_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_123_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16461_ clknet_leaf_21_wb_clk_i _02215_ _00444_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13673_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[28\] net567 net345 team_01_WB.instance_to_wrap.cpu.f0.i\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10885_ net516 _07041_ _07099_ _07224_ vssd1 vssd1 vccd1 vccd1 _07225_ sky130_fd_sc_hd__a31o_1
XANTENNA__11660__X _07866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15412_ net1379 vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12624_ net2717 net218 net392 vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__mux2_1
X_16392_ clknet_leaf_95_wb_clk_i net2533 _00375_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[115\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17995__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15343_ net1391 vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12555_ _07942_ _07951_ net573 vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__and3_4
XANTENNA__12408__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11506_ net1810 net877 _07758_ _07780_ vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__o22a_1
X_15274_ net1295 vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__inv_2
X_12486_ net2296 net319 net414 vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17013_ clknet_leaf_114_wb_clk_i _02700_ _00996_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14225_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[7\] vssd1 vssd1 vccd1
+ vccd1 _02262_ sky130_fd_sc_hd__clkbuf_1
X_11437_ net1070 _07700_ net324 vssd1 vssd1 vccd1 vccd1 _07743_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08397__A1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14156_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[1\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11368_ _07696_ vssd1 vssd1 vccd1 vccd1 _07697_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13107_ net73 net71 net74 _03729_ vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__and4_1
XANTENNA__12143__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10319_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[18\] net787 net742 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[18\]
+ _06658_ vssd1 vssd1 vccd1 vccd1 _06659_ sky130_fd_sc_hd__a221o_1
XANTENNA__10452__A net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14087_ _04365_ _04374_ vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__or2_1
X_11299_ net197 net193 net643 vssd1 vssd1 vccd1 vccd1 _07639_ sky130_fd_sc_hd__o21ai_4
XANTENNA__09346__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17915_ net1522 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
X_13038_ net2897 net2832 net857 vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__mux2_1
XANTENNA__14859__A net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11982__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1150 net1151 vssd1 vssd1 vccd1 vccd1 net1150 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13763__A net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1161 net1163 vssd1 vssd1 vccd1 vccd1 net1161 sky130_fd_sc_hd__clkbuf_2
Xfanout1172 team_01_WB.instance_to_wrap.cpu.DM0.ihit vssd1 vssd1 vccd1 vccd1 net1172
+ sky130_fd_sc_hd__clkbuf_2
X_17846_ clknet_leaf_120_wb_clk_i _03522_ _01786_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[116\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout1183 net1185 vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08857__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1194 net1201 vssd1 vssd1 vccd1 vccd1 net1194 sky130_fd_sc_hd__buf_2
XFILLER_0_89_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14989_ net1265 vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__inv_2
X_17777_ clknet_leaf_121_wb_clk_i net2775 _01717_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16728_ clknet_leaf_49_wb_clk_i _02415_ _00711_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16659_ clknet_leaf_18_wb_clk_i _02346_ _00642_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08872__A2 _04806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09200_ net1082 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[17\] net892
+ vssd1 vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__and3_1
XANTENNA__11208__A1 _06920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_971 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12956__A1 _05110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09131_ net1022 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[14\] net937 vssd1
+ vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12318__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08624__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09062_ net1029 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[12\] net902
+ vssd1 vssd1 vccd1 vccd1 _05402_ sky130_fd_sc_hd__and3_1
XANTENNA_wire583_X net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire962_A _04656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10431__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_96_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08013_ net1427 vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold600 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2135 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold611 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[15\] vssd1 vssd1 vccd1 vccd1
+ net2146 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_25_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_130_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold622 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2168 sky130_fd_sc_hd__dlygate4sd3_1
Xhold644 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2179 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold655 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2190 sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[26\] vssd1 vssd1 vccd1 vccd1
+ net2212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 _02089_ vssd1 vssd1 vccd1 vccd1 net2223 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12053__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold699 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2234 sky130_fd_sc_hd__dlygate4sd3_1
X_09964_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[3\] net816 net802 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[3\]
+ _06299_ vssd1 vssd1 vccd1 vccd1 _06304_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1115_A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08915_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[2\] net651 _05227_ _05244_
+ _05247_ vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_55_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13944__Y _04236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09895_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[5\] net820 net757 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06235_ sky130_fd_sc_hd__a22o_1
Xhold1300 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2835 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1311 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[30\] vssd1 vssd1 vccd1 vccd1
+ net2846 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1322 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2857 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_86_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08846_ _05160_ _05183_ _05184_ _05185_ vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__or4_1
Xhold1333 team_01_WB.instance_to_wrap.cpu.c0.count\[4\] vssd1 vssd1 vccd1 vccd1 net2868
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1344 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1355 team_01_WB.instance_to_wrap.cpu.c0.count\[8\] vssd1 vssd1 vccd1 vccd1 net2890
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1366 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2901 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1377 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[78\] vssd1 vssd1 vccd1 vccd1
+ net2912 sky130_fd_sc_hd__dlygate4sd3_1
X_08777_ net1093 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[0\] net905 vssd1
+ vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout742_A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1388 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2923 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout363_X net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13960__X _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1399 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2934 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_0_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11447__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10655__C1 _05263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout530_X net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout628_X net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10670_ net552 _06398_ vssd1 vssd1 vccd1 vccd1 _07010_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08933__C net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08076__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09329_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[24\] net691 net687 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[24\]
+ _05668_ vssd1 vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__a221o_1
XANTENNA__10096__X _06436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12228__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08615__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14149__B1 _04266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12340_ net2548 net263 net427 vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08007__A net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout997_X net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12271_ net3080 net239 net435 vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_33_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14010_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[73\] _04235_ _04255_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[113\]
+ _04294_ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__a221o_1
X_11222_ net556 _06980_ _07132_ _07560_ _07561_ vssd1 vssd1 vccd1 vccd1 _07562_ sky130_fd_sc_hd__o311ai_1
XANTENNA__13372__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10186__A1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11368__A _07696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11153_ _06254_ _06255_ _06284_ _06409_ vssd1 vssd1 vccd1 vccd1 _07493_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_105_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_147_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09328__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10104_ net1156 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[6\] net964 vssd1
+ vssd1 vccd1 vccd1 _06444_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11084_ _05729_ _06811_ _07344_ vssd1 vssd1 vccd1 vccd1 _07424_ sky130_fd_sc_hd__or3b_1
X_15961_ net1403 vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__inv_2
XANTENNA__14679__A net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1071 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10035_ net1142 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[0\] net957 vssd1
+ vssd1 vccd1 vccd1 _06375_ sky130_fd_sc_hd__and3_1
XANTENNA__11655__X _07862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17700_ clknet_leaf_137_wb_clk_i _03384_ _01641_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[21\]
+ sky130_fd_sc_hd__dfrtp_4
X_14912_ net1235 vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_125_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11686__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15892_ net1360 vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__inv_2
XANTENNA__08677__A net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17631_ clknet_leaf_3_wb_clk_i _03316_ _01572_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14843_ net1254 vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17562_ clknet_leaf_89_wb_clk_i _03249_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_14774_ net1253 vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__inv_2
X_11986_ net2535 net292 net474 vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__mux2_1
X_16513_ clknet_leaf_5_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[11\]
+ _00496_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16920__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13725_ _04109_ _04131_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[14\]
+ sky130_fd_sc_hd__nor2_1
X_10937_ _07067_ _07157_ net514 vssd1 vssd1 vccd1 vccd1 _07277_ sky130_fd_sc_hd__mux2_1
X_17493_ clknet_leaf_114_wb_clk_i _03180_ _01476_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09004__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12927__A net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16444_ clknet_leaf_42_wb_clk_i _02198_ _00427_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13656_ _03872_ _03876_ vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__xor2_1
X_10868_ _06740_ _07112_ _06715_ vssd1 vssd1 vccd1 vccd1 _07208_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_72_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_94_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12607_ net3123 net254 net396 vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__mux2_1
XANTENNA__12938__B2 net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16375_ clknet_leaf_90_wb_clk_i net2899 _00358_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[98\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13587_ _03902_ _04031_ vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12138__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10799_ _07137_ _07138_ net519 vssd1 vssd1 vccd1 vccd1 _07139_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15326_ net1316 vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__inv_2
X_12538_ net2184 net263 net404 vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11977__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15257_ net1233 vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12469_ net2915 net238 net411 vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__mux2_1
X_14208_ net2326 vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__clkbuf_1
X_17891__1513 vssd1 vssd1 vccd1 vccd1 net1513 _17891__1513/LO sky130_fd_sc_hd__conb_1
XANTENNA__09674__C net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15188_ net1379 vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__inv_2
XANTENNA__09031__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14139_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[95\] _04240_ _04250_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[127\]
+ _04423_ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout409 _03564_ vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_33_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08700_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[7\] net702 _05036_ _05039_
+ vssd1 vssd1 vccd1 vccd1 _05040_ sky130_fd_sc_hd__o22ai_4
XANTENNA__12601__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09680_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[22\] net794 _06010_ _06012_
+ _06013_ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12874__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08448__A_N net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08587__A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08542__A1 net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_143_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_143_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08631_ team_01_WB.instance_to_wrap.cpu.CU0.bit30 net596 vssd1 vssd1 vccd1 vccd1
+ _04971_ sky130_fd_sc_hd__nand2_2
X_17829_ clknet_leaf_96_wb_clk_i net2237 _01769_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[99\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08562_ net1078 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[19\] net922
+ vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_81_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14091__A2 _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17949__1464 vssd1 vssd1 vccd1 vccd1 _17949__1464/HI net1464 sky130_fd_sc_hd__conb_1
XANTENNA__10637__C1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08493_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[23\] net676 _04809_
+ _04824_ _04769_ vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_9_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08845__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08753__C net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09211__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12048__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout323_A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1065_A team_01_WB.instance_to_wrap.cpu.RU0.state\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09114_ _05418_ net584 net601 vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__mux2_2
XFILLER_0_5_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11887__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09045_ net1110 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[12\] net924
+ vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1232_A net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09558__B1 _05897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11459__Y _07755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold430 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1965 sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1976 sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1987 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout692_A net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold463 team_01_WB.instance_to_wrap.a1.ADR_I\[8\] vssd1 vssd1 vccd1 vccd1 net1998
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13955__X _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold474 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2009 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1020_X net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold485 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2020 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1118_X net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_117_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold496 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2031 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10523__C net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout910 net913 vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__buf_4
X_09947_ net1155 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[3\] _04640_
+ vssd1 vssd1 vccd1 vccd1 _06287_ sky130_fd_sc_hd__and3_1
Xfanout932 net933 vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout480_X net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout943 net944 vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__clkbuf_8
Xfanout954 net955 vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__buf_4
XFILLER_0_99_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout578_X net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout965 _04650_ vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__buf_4
XANTENNA__12511__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout976 _04638_ vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__buf_4
Xfanout987 net989 vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__clkbuf_4
X_09878_ _06217_ net341 vssd1 vssd1 vccd1 vccd1 _06218_ sky130_fd_sc_hd__nand2b_2
XTAP_TAPCELL_ROW_70_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1130 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2665 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout998 _04491_ vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__clkbuf_4
Xhold1141 _03479_ vssd1 vssd1 vccd1 vccd1 net2676 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08928__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08829_ net1022 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[1\] net907 vssd1
+ vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__and3_1
Xhold1152 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[46\] vssd1 vssd1 vccd1 vccd1
+ net2687 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1163 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2698 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout745_X net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1174 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[119\] vssd1 vssd1 vccd1 vccd1
+ net2709 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1185 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 net2720
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1196 _03500_ vssd1 vssd1 vccd1 vccd1 net2731 sky130_fd_sc_hd__dlygate4sd3_1
X_11840_ net1840 net233 net487 vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14082__A2 _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout912_X net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11771_ net2292 net238 net495 vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__mux2_1
XANTENNA__08836__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13847__A_N net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13510_ _03844_ _03948_ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10722_ net534 _07010_ vssd1 vssd1 vccd1 vccd1 _07062_ sky130_fd_sc_hd__or2_2
X_14490_ net1356 vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13441_ _05456_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] vssd1 vssd1
+ vccd1 vccd1 _03902_ sky130_fd_sc_hd__and2b_1
X_10653_ _04706_ net543 net536 _06992_ vssd1 vssd1 vccd1 vccd1 _06993_ sky130_fd_sc_hd__o211a_1
XANTENNA__10267__A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16160_ clknet_leaf_131_wb_clk_i _01923_ _00148_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12871__A_N net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08382__D _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13372_ net1567 net829 _03838_ team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1
+ vccd1 vccd1 _01875_ sky130_fd_sc_hd__a22o_1
X_10584_ _06901_ _06917_ vssd1 vssd1 vccd1 vccd1 _06924_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_118_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09261__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload19 clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload19/Y sky130_fd_sc_hd__inv_6
X_15111_ net1389 vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_118_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_156_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11797__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12323_ net2437 net290 net432 vssd1 vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__mux2_1
X_16091_ clknet_leaf_132_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[13\]
+ _00079_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[13\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09549__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15042_ net1320 vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__inv_2
X_12254_ net2744 net305 net442 vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__mux2_1
XANTENNA__10714__B _06928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13728__D _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11205_ net373 net334 net332 vssd1 vssd1 vccd1 vccd1 _07545_ sky130_fd_sc_hd__a21o_1
X_12185_ net2277 net310 net447 vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11136_ _07469_ _07470_ _07475_ vssd1 vssd1 vccd1 vccd1 _07476_ sky130_fd_sc_hd__a21bo_2
XANTENNA__08772__B2 net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16993_ clknet_leaf_55_wb_clk_i _02680_ _00976_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11067_ _07368_ _07405_ _04947_ net374 vssd1 vssd1 vccd1 vccd1 _07407_ sky130_fd_sc_hd__o2bb2a_1
X_15944_ net1402 vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__inv_2
XANTENNA__12421__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10018_ _06346_ _06349_ _06354_ _06357_ vssd1 vssd1 vccd1 vccd1 _06358_ sky130_fd_sc_hd__or4_1
X_15875_ net1309 vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14826_ net1374 vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__inv_2
X_17614_ clknet_leaf_2_wb_clk_i _03299_ _01555_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14073__A2 _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17545_ clknet_leaf_40_wb_clk_i _03232_ _01528_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14757_ net1274 vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__inv_2
X_11969_ net2199 net202 net472 vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13105__X net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13708_ team_01_WB.instance_to_wrap.cpu.c0.count\[1\] team_01_WB.instance_to_wrap.cpu.c0.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__or2_1
X_17476_ clknet_leaf_82_wb_clk_i _03163_ _01459_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_14688_ net1204 vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09669__C net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08573__C net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16427_ clknet_leaf_140_wb_clk_i _02181_ _00410_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13639_ net725 _07308_ net987 vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14872__A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16358_ clknet_leaf_87_wb_clk_i _02112_ _00341_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[81\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10398__A1 _06737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09252__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15309_ net1265 vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16289_ clknet_leaf_118_wb_clk_i _02043_ _00272_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[12\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_140_832 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_11__f_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout206 net209 vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__buf_2
X_09801_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[14\] net800 _06139_
+ _06140_ vssd1 vssd1 vccd1 vccd1 _06141_ sky130_fd_sc_hd__a211o_1
XANTENNA__10343__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout217 _07835_ vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09960__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout228 _07900_ vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__buf_2
XANTENNA__13935__B team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07993_ net1137 vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__inv_2
Xfanout239 net240 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__buf_2
XFILLER_0_66_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13639__A2 _07308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09732_ net1145 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[20\] net982
+ vssd1 vssd1 vccd1 vccd1 _06072_ sky130_fd_sc_hd__and3_1
XANTENNA__12331__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08748__C _04779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09663_ net1144 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[22\] net980
+ vssd1 vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__and3_1
XANTENNA__08110__A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08614_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[11\] net690 net672 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_19_Left_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09594_ net512 _05933_ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14064__A2 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08279__A0 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08545_ net1134 net620 net593 vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout440_A _07962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout538_A net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08476_ net1001 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[23\] net878
+ vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_46_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09491__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout705_A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout326_X net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_40_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_31_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire618 _05331_ vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__clkbuf_1
XANTENNA__13575__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09779__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09243__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08987__D1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13398__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_28_Left_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12506__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1235_X net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13327__A1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09028_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[9\] net679 _05340_ _05350_
+ _05361_ vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_142_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout695_X net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold260 _01996_ vssd1 vssd1 vccd1 vccd1 net1795 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10026__S _04628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold271 _03310_ vssd1 vssd1 vccd1 vccd1 net1806 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_72_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold282 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[2\] vssd1 vssd1 vccd1 vccd1
+ net1817 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10010__B1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold293 team_01_WB.instance_to_wrap.a1.ADR_I\[6\] vssd1 vssd1 vccd1 vccd1 net1828
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout740 net741 vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_1053 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout751 net752 vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__clkbuf_8
Xfanout762 _04674_ vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12241__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13990_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[112\] _04255_ _04260_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[56\]
+ _04272_ vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__a221o_1
Xfanout773 net774 vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout784 _04661_ vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__clkbuf_8
Xfanout795 net797 vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11365__B team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12941_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[10\] net1038 vssd1 vssd1 vccd1
+ vccd1 _03704_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_37_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10959__A1_N _06958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15660_ net1259 vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__inv_2
X_12872_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[31\] _03654_ net1040 vssd1
+ vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__mux2_1
X_14611_ net1323 vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__inv_2
X_11823_ net2100 net288 net492 vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__mux2_1
X_15591_ net1395 vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__inv_2
XANTENNA__13263__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_96_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13072__S net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17330_ clknet_leaf_145_wb_clk_i _03017_ _01313_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_14542_ net1354 vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__inv_2
X_11754_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[0\] _07438_ net715 vssd1 vssd1
+ vccd1 vccd1 _07940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_7__f_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10705_ _05805_ net513 vssd1 vssd1 vccd1 vccd1 _07045_ sky130_fd_sc_hd__xor2_2
X_17261_ clknet_leaf_108_wb_clk_i _02948_ _01244_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_14473_ net1358 vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__inv_2
X_11685_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[14\] net713 vssd1 vssd1 vccd1
+ vccd1 _07885_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16212_ clknet_leaf_124_wb_clk_i net1923 _00200_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13566__A1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13424_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] _04949_ _03884_ vssd1
+ vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__nor3_1
XANTENNA__09786__A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17192_ clknet_leaf_62_wb_clk_i _02879_ _01175_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10636_ _06912_ _06919_ _06975_ vssd1 vssd1 vccd1 vccd1 _06976_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09234__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload108 clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload108/Y sky130_fd_sc_hd__clkinv_8
X_16143_ clknet_leaf_137_wb_clk_i _01906_ _00131_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload119 clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload119/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_106_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13355_ team_01_WB.instance_to_wrap.cpu.f0.i\[9\] net1070 team_01_WB.instance_to_wrap.cpu.f0.i\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12416__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10567_ net512 net511 net543 vssd1 vssd1 vccd1 vccd1 _06907_ sky130_fd_sc_hd__mux2_1
X_12306_ net2692 net267 net432 vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__mux2_1
X_16074_ clknet_leaf_153_wb_clk_i _01867_ _00062_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\]
+ sky130_fd_sc_hd__dfstp_4
XFILLER_0_122_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13286_ _03773_ _03771_ net825 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[27\]
+ vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__o2bb2a_1
X_10498_ net1131 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[31\] net948
+ vssd1 vssd1 vccd1 vccd1 _06838_ sky130_fd_sc_hd__and3_1
X_15025_ net1393 vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__inv_2
X_17948__1463 vssd1 vssd1 vccd1 vccd1 _17948__1463/HI net1463 sky130_fd_sc_hd__conb_1
X_12237_ net3016 net269 net439 vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__mux2_1
XANTENNA__10001__B1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12168_ net2216 net241 net449 vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__mux2_1
XANTENNA__09952__C net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10552__A1 _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11119_ net558 _07456_ _07458_ vssd1 vssd1 vccd1 vccd1 _07459_ sky130_fd_sc_hd__o21a_1
XANTENNA__12151__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12829__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16976_ clknet_leaf_145_wb_clk_i _02663_ _00959_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_12099_ net2397 net273 net457 vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__mux2_1
Xinput6 DAT_I[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_3_4_0_wb_clk_i_X clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15927_ net1413 vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__inv_2
XANTENNA__11990__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15858_ net1356 vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__inv_2
XANTENNA__08865__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14046__A2 _04221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1060 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_wire506_A _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14809_ net1238 vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15789_ net1191 vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__inv_2
X_08330_ net995 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[30\] net956 vssd1
+ vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__and3_1
X_17528_ clknet_leaf_38_wb_clk_i _03215_ _01511_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08261_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[20\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[12\]
+ net1045 vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17459_ clknet_leaf_20_wb_clk_i _03146_ _01442_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10338__C net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08192_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[89\] net2799 net1057 vssd1 vssd1
+ vccd1 vccd1 _03495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16590__Q team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[22\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12326__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10240__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10791__B2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10073__C net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1028_A net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08736__A1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09933__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout390_A _03569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout488_A _07947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10370__A net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12061__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07976_ team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1 _04474_
+ sky130_fd_sc_hd__inv_2
X_09715_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[21\] net746 _06041_ _06042_
+ _06048_ vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08478__C net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12296__A1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout655_A _04817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1397_A net1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09646_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[23\] net730 _05969_ _05973_
+ _05975_ vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__a2111o_1
XANTENNA__14037__A2 _04265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[25\] net812 net773 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout822_A net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout443_X net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1185_X net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08528_ net1077 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[18\] net918
+ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_65_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08459_ net1116 net1119 net1122 net1125 vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__and4bb_4
XANTENNA__09102__C net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout708_X net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13548__A1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11470_ net366 _07762_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[28\] net874
+ vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09216__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_154_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08941__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10421_ net1133 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[27\] net975
+ vssd1 vssd1 vccd1 vccd1 _06761_ sky130_fd_sc_hd__and3b_1
XFILLER_0_150_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12236__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10231__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12771__A2 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13140_ net1686 net846 net634 team_01_WB.instance_to_wrap.a1.ADR_I\[3\] vssd1 vssd1
+ vccd1 vccd1 _02001_ sky130_fd_sc_hd__a22o_1
X_10352_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[17\] net736 net733 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _06692_ sky130_fd_sc_hd__a22o_1
XANTENNA__08015__A _04504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13071_ net2883 net2854 net856 vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11079__C _05657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10283_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[19\] net776 net759 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _06623_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12022_ net2396 net317 net469 vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__mux2_1
XANTENNA_input49_A wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_10__f_wb_clk_i_X clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16830_ clknet_leaf_80_wb_clk_i _02517_ _00813_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_45_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout570 _04520_ vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__buf_2
XANTENNA__17637__CLK clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16761_ clknet_leaf_102_wb_clk_i _02448_ _00744_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13973_ _04217_ _04222_ _04239_ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_109_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12924_ _04944_ _07752_ net361 vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__a21oi_4
X_15712_ net1242 vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__inv_2
X_16692_ clknet_leaf_66_wb_clk_i _02379_ _00675_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14028__A2 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12919__B net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12039__A1 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12855_ net2849 net251 net381 vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__mux2_1
X_15643_ net1251 vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__inv_2
X_11806_ net2962 net265 net492 vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__mux2_1
X_15574_ net1261 vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12786_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[14\] net304 net1037 vssd1 vssd1
+ vccd1 vccd1 _03619_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09455__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17313_ clknet_leaf_54_wb_clk_i _03000_ _01296_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_14525_ net1412 vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__inv_2
X_11737_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[4\] net716 vssd1 vssd1 vccd1
+ vccd1 _07927_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_54_Left_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09012__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10470__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17244_ clknet_leaf_58_wb_clk_i _02931_ _01227_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_14456_ net1224 vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__inv_2
X_11668_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] _07812_ vssd1 vssd1
+ vccd1 vccd1 _07872_ sky130_fd_sc_hd__xor2_1
XFILLER_0_22_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09947__C _04640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08851__C net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13407_ _03866_ _03867_ vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10619_ _06945_ _06958_ net528 vssd1 vssd1 vccd1 vccd1 _06959_ sky130_fd_sc_hd__mux2_1
X_17175_ clknet_leaf_14_wb_clk_i _02862_ _01158_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12146__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14387_ net1186 vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwire960 net961 vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__clkbuf_2
X_11599_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] _07814_ vssd1 vssd1
+ vccd1 vccd1 _07816_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_12_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10222__B1 _06560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16126_ clknet_leaf_126_wb_clk_i _00007_ _00114_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__12762__A2 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13338_ _07682_ _03812_ _03813_ vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_40_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11985__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16057_ clknet_leaf_4_wb_clk_i _01850_ _00045_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\]
+ sky130_fd_sc_hd__dfrtp_4
X_13269_ team_01_WB.instance_to_wrap.cpu.f0.i\[28\] net1068 _03754_ _03755_ net564
+ vssd1 vssd1 vccd1 vccd1 _03760_ sky130_fd_sc_hd__o311a_1
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15008_ net1235 vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_63_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11722__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11286__A _07019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10190__A _06526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16959_ clknet_leaf_44_wb_clk_i _02646_ _00942_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_09500_ net997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[29\] net949 vssd1
+ vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__and3_1
XANTENNA__14019__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16585__Q team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[17\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09431_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[28\] net691 net687 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[28\]
+ _05770_ vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09362_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[25\] _04766_ net655
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[25\] _05701_ vssd1 vssd1 vccd1
+ vccd1 _05702_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_23_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08313_ net1158 net1161 net1164 net1166 vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__and4b_2
XTAP_TAPCELL_ROW_43_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09293_ net1003 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[22\] net918 vssd1
+ vssd1 vccd1 vccd1 _05633_ sky130_fd_sc_hd__and3_1
XANTENNA_11 _03663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout236_A _07873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_33 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08244_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[37\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[29\]
+ net1051 vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__mux2_1
XANTENNA_44 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09857__C net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_55 _03654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_66 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08175_ net2943 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[98\] net1052 vssd1 vssd1
+ vccd1 vccd1 _03512_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12056__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10365__A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout403_A net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_6__f_wb_clk_i_X clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1145_A net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10213__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12753__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10764__A1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11895__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput140 net140 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1312_A net1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput151 net151 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
Xoutput162 net162 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__clkbuf_4
XANTENNA__09906__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput173 net173 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__clkbuf_4
Xoutput184 net184 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout772_A net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout393_X net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13963__X _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout560_X net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout658_X net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10970_ _06255_ _06410_ _07291_ _07309_ net344 vssd1 vssd1 vccd1 vccd1 _07310_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_67_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09685__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08936__C net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09629_ net1135 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[23\] net963
+ vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_104_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12640_ net1987 net255 net394 vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__mux2_1
X_17947__1462 vssd1 vssd1 vccd1 vccd1 _17947__1462/HI net1462 sky130_fd_sc_hd__conb_1
XANTENNA__09437__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_156_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12571_ net2156 net264 net400 vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_156_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12755__A net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14310_ net1324 vssd1 vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11522_ net2276 net1171 net588 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1
+ vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15290_ net1313 vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08671__C net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14241_ net1229 vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__inv_2
X_11453_ net1175 _04621_ _07669_ team_01_WB.instance_to_wrap.cpu.f0.i\[0\] vssd1 vssd1
+ vccd1 vccd1 _07751_ sky130_fd_sc_hd__a31o_1
XFILLER_0_135_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10275__A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10404_ _06598_ _06604_ _06743_ vssd1 vssd1 vccd1 vccd1 _06744_ sky130_fd_sc_hd__a21o_1
X_14172_ net1426 _04446_ _04447_ vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__nor3_1
XFILLER_0_21_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11384_ team_01_WB.instance_to_wrap.cpu.f0.i\[23\] _07712_ vssd1 vssd1 vccd1 vccd1
+ _07713_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13123_ net1735 net843 net631 team_01_WB.instance_to_wrap.a1.ADR_I\[20\] vssd1 vssd1
+ vccd1 vccd1 _02018_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10335_ _06673_ _06674_ _06672_ vssd1 vssd1 vccd1 vccd1 _06675_ sky130_fd_sc_hd__a21o_1
XANTENNA__10562__X _06902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17931_ net1448 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
X_13054_ net2637 net2388 net857 vssd1 vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__mux2_1
X_10266_ net1128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[19\] net965
+ vssd1 vssd1 vccd1 vccd1 _06606_ sky130_fd_sc_hd__and3_1
Xfanout1310 net1322 vssd1 vssd1 vccd1 vccd1 net1310 sky130_fd_sc_hd__clkbuf_2
X_12005_ net1883 net237 net467 vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__mux2_1
Xfanout1321 net1322 vssd1 vssd1 vccd1 vccd1 net1321 sky130_fd_sc_hd__clkbuf_4
Xfanout1332 net1430 vssd1 vssd1 vccd1 vccd1 net1332 sky130_fd_sc_hd__clkbuf_2
X_17862_ clknet_leaf_125_wb_clk_i _03537_ _01802_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10197_ net1140 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[8\] net965 vssd1
+ vssd1 vccd1 vccd1 _06537_ sky130_fd_sc_hd__and3_1
Xfanout1343 net1344 vssd1 vssd1 vccd1 vccd1 net1343 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11180__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1354 net1355 vssd1 vssd1 vccd1 vccd1 net1354 sky130_fd_sc_hd__buf_4
Xfanout1365 net1369 vssd1 vssd1 vccd1 vccd1 net1365 sky130_fd_sc_hd__buf_2
X_16813_ clknet_leaf_108_wb_clk_i _02500_ _00796_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_128_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1376 net1377 vssd1 vssd1 vccd1 vccd1 net1376 sky130_fd_sc_hd__buf_2
XFILLER_0_75_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09007__C net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1387 net1398 vssd1 vssd1 vccd1 vccd1 net1387 sky130_fd_sc_hd__buf_4
XANTENNA__12489__X _03564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17793_ clknet_leaf_122_wb_clk_i _03469_ _01733_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[63\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1398 net1429 vssd1 vssd1 vccd1 vccd1 net1398 sky130_fd_sc_hd__buf_4
X_16744_ clknet_leaf_60_wb_clk_i _02431_ _00727_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13956_ _04223_ _04231_ vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__nand2_2
XANTENNA__09676__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12907_ _05615_ net578 net361 vssd1 vssd1 vccd1 vccd1 _03680_ sky130_fd_sc_hd__o21ba_1
X_13887_ _04193_ vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__inv_2
X_16675_ clknet_leaf_26_wb_clk_i _02362_ _00658_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_12838_ net2376 net210 net379 vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__mux2_1
X_15626_ net1374 vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09428__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15557_ net1288 vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__inv_2
X_12769_ net1966 net638 net606 _03607_ vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14508_ net1407 vssd1 vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15488_ net1270 vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08581__C net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput20 DAT_I[26] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
X_17227_ clknet_leaf_9_wb_clk_i _02914_ _01210_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_14439_ net1306 vssd1 vssd1 vccd1 vccd1 _00233_ sky130_fd_sc_hd__inv_2
Xinput31 DAT_I[7] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput42 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_1
Xinput53 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_1
Xinput64 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_25_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17158_ clknet_leaf_90_wb_clk_i _02845_ _01141_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16557__CLK clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold804 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2339 sky130_fd_sc_hd__dlygate4sd3_1
Xhold815 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[114\] vssd1 vssd1 vccd1 vccd1
+ net2350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09600__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold826 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold837 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[42\] vssd1 vssd1 vccd1 vccd1
+ net2372 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10746__B2 _05263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16109_ clknet_leaf_138_wb_clk_i _01884_ _00097_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold848 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2383 sky130_fd_sc_hd__dlygate4sd3_1
X_17089_ clknet_leaf_55_wb_clk_i _02776_ _01072_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_09980_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[2\] net818 net773 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[2\]
+ _06319_ vssd1 vssd1 vccd1 vccd1 _06320_ sky130_fd_sc_hd__a221o_1
XANTENNA__12604__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold859 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2394 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08931_ net1107 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[6\] net915 vssd1
+ vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13160__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08862_ net1106 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[3\] net898 vssd1
+ vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_36_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1504 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net3039 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1515 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net3050 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1526 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net3061 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_88_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08793_ _05120_ _05124_ _05128_ _05132_ vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__or4_1
Xhold1537 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net3072 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_88_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1548 team_01_WB.instance_to_wrap.cpu.K0.code\[4\] vssd1 vssd1 vccd1 vccd1 net3083
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09116__A1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold1559 team_01_WB.instance_to_wrap.cpu.K0.code\[7\] vssd1 vssd1 vccd1 vccd1 net3094
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout186_A _07639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08756__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1095_A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10682__A0 _04706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09414_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[27\] net693 net674 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[27\]
+ _05740_ vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09345_ net1115 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[25\] net942
+ vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout520_A _05260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10434__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09276_ net1127 net711 net594 vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__a21o_1
XFILLER_0_106_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15886__A net1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08227_ net2737 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[46\] net1043 vssd1 vssd1
+ vccd1 vccd1 _03460_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_151_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout406_X net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1148_X net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09884__A net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08158_ net1782 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[115\] net1054 vssd1 vssd1
+ vccd1 vccd1 _03529_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout987_A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12514__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08089_ _04523_ _04530_ _04536_ _04542_ vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__or4_1
X_10120_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[6\] net788 _04667_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[6\]
+ _06459_ vssd1 vssd1 vccd1 vccd1 _06460_ sky130_fd_sc_hd__a221o_1
XANTENNA__11638__B _07600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout775_X net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10051_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[0\] net804 net790 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06391_ sky130_fd_sc_hd__a22o_1
XANTENNA__13151__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout942_X net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13853__B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11654__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13810_ net2664 net833 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[3\]
+ sky130_fd_sc_hd__and2_1
X_14790_ net1381 vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__inv_2
XANTENNA__09124__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13741_ net1178 net2195 net1061 vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__a21o_1
X_10953_ _06441_ _06470_ vssd1 vssd1 vccd1 vccd1 _07293_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_123_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_123_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13672_ net1628 net568 net347 team_01_WB.instance_to_wrap.cpu.f0.i\[29\] vssd1 vssd1
+ vccd1 vccd1 _01830_ sky130_fd_sc_hd__a22o_1
X_16460_ clknet_leaf_28_wb_clk_i _02214_ _00443_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10884_ net333 _07222_ _07223_ net336 vssd1 vssd1 vccd1 vccd1 _07224_ sky130_fd_sc_hd__a22o_1
XANTENNA__08963__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15411_ net1394 vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__inv_2
X_12623_ net2417 net224 net391 vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__mux2_1
X_16391_ clknet_leaf_88_wb_clk_i _02145_ _00374_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[114\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_62_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08618__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13080__S net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15342_ net1300 vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10425__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12554_ net1778 net291 net406 vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__mux2_1
XANTENNA__12965__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10976__A1 _07015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09830__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11505_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[10\] _07756_ vssd1 vssd1 vccd1
+ vccd1 _07780_ sky130_fd_sc_hd__and2_1
X_15273_ net1293 vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__inv_2
X_12485_ net2182 net307 net414 vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14224_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[8\] vssd1 vssd1 vccd1
+ vccd1 _02263_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_input71_X net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09794__A net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17012_ clknet_leaf_21_wb_clk_i _02699_ _00995_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11436_ team_01_WB.instance_to_wrap.cpu.f0.i\[9\] _07736_ _07742_ vssd1 vssd1 vccd1
+ vccd1 _03372_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_145_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12932__B net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14155_ net1696 _04195_ net1421 vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_145_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11367_ _04575_ _07651_ vssd1 vssd1 vccd1 vccd1 _07696_ sky130_fd_sc_hd__or2_2
XANTENNA__12424__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13106_ net179 vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10318_ net990 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[18\] net945 vssd1
+ vssd1 vccd1 vccd1 _06658_ sky130_fd_sc_hd__o21a_1
X_14086_ _04367_ _04369_ _04371_ _04373_ vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__or4_1
X_11298_ net1075 _07637_ vssd1 vssd1 vccd1 vccd1 _07638_ sky130_fd_sc_hd__nand2_1
X_13037_ net2444 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[57\] net865 vssd1 vssd1
+ vccd1 vccd1 _02088_ sky130_fd_sc_hd__mux2_1
XANTENNA__13142__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17914_ net1445 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
X_10249_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[9\] net767 _06583_ _06588_
+ vssd1 vssd1 vccd1 vccd1 _06589_ sky130_fd_sc_hd__o22a_2
Xfanout1140 net1141 vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__buf_1
XANTENNA__09897__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1151 net1157 vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__clkbuf_2
Xfanout1162 net1163 vssd1 vssd1 vccd1 vccd1 net1162 sky130_fd_sc_hd__clkbuf_2
X_17845_ clknet_leaf_96_wb_clk_i net1749 _01785_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[115\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10900__A1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1173 net1174 vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__buf_2
Xfanout1184 net1185 vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__clkbuf_2
Xfanout1195 net1201 vssd1 vssd1 vccd1 vccd1 net1195 sky130_fd_sc_hd__buf_4
XFILLER_0_89_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17776_ clknet_leaf_117_wb_clk_i net2586 _01716_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[46\]
+ sky130_fd_sc_hd__dfrtp_1
X_14988_ net1260 vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09649__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11283__B _07232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16727_ clknet_leaf_15_wb_clk_i _02414_ _00710_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13939_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__nor2_2
XFILLER_0_88_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16658_ clknet_leaf_144_wb_clk_i _02345_ _00641_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15609_ net1237 vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08609__B1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13602__B1 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16589_ clknet_leaf_144_wb_clk_i _02276_ _00572_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[21\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_151_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09130_ net1024 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[14\] net919 vssd1
+ vssd1 vccd1 vccd1 _05470_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09040__Y _05380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10186__Y _06526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10627__B net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10967__A1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09061_ net1109 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[12\] net915
+ vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__and3_1
XANTENNA__09200__C net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10346__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08012_ net1 vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__inv_2
Xhold601 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2136 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold612 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2147 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold623 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1 net2158
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold634 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2169 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12334__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap342 _05378_ vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_38_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold645 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2180 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold656 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold667 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[16\] vssd1 vssd1 vccd1 vccd1
+ net2202 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_107_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09209__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09963_ _06286_ _06300_ _06301_ _06302_ vssd1 vssd1 vccd1 vccd1 _06303_ sky130_fd_sc_hd__or4_1
Xhold678 _03440_ vssd1 vssd1 vccd1 vccd1 net2213 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13669__A0 net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold689 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[10\] vssd1 vssd1 vccd1 vccd1
+ net2224 sky130_fd_sc_hd__dlygate4sd3_1
X_17946__1461 vssd1 vssd1 vccd1 vccd1 _17946__1461/HI net1461 sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_65_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08914_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[2\] net659 _05243_ _05245_
+ net707 vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13133__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16103__Q team_01_WB.instance_to_wrap.cpu.f0.data_adr\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1010_A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09894_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[5\] net800 net783 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06234_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1108_A net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1301 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[47\] vssd1 vssd1 vccd1 vccd1
+ net2836 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1312 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[11\] vssd1 vssd1 vccd1 vccd1
+ net2847 sky130_fd_sc_hd__dlygate4sd3_1
X_08845_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[1\] net662 net657 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__a22o_1
Xhold1323 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[102\] vssd1 vssd1 vccd1 vccd1
+ net2858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1334 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1345 team_01_WB.instance_to_wrap.cpu.K0.enable vssd1 vssd1 vccd1 vccd1 net2880
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1356 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2891 sky130_fd_sc_hd__dlygate4sd3_1
X_08776_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] _04751_ _04752_ net1127 vssd1
+ vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__a22o_4
Xhold1367 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2902 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1378 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2913 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14094__B1 _04266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1389 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2924 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08486__C net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11193__B net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout356_X net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout735_A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1098_X net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout902_A net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12509__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09328_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[24\] net699 net655 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__a22o_1
XANTENNA__09273__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09812__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11080__B1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09259_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[20\] net680 net676 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[20\]
+ _05596_ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_146_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_90_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09818__S _04628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12270_ net2965 net270 net435 vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__mux2_1
XANTENNA__13848__B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout892_X net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11221_ net556 _07202_ _07017_ vssd1 vssd1 vccd1 vccd1 _07561_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12244__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10186__A2 _06525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11152_ _06284_ _06409_ _06254_ _06255_ vssd1 vssd1 vccd1 vccd1 _07492_ sky130_fd_sc_hd__o211a_1
X_10103_ net1155 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[6\] net985 vssd1
+ vssd1 vccd1 vccd1 _06443_ sky130_fd_sc_hd__and3_1
XANTENNA__13124__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11083_ _05681_ net511 _07349_ _05707_ net512 vssd1 vssd1 vccd1 vccd1 _07423_ sky130_fd_sc_hd__o32a_1
X_15960_ net1354 vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__inv_2
XANTENNA__11135__B2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input31_A DAT_I[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10034_ net1142 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[0\] net954 vssd1
+ vssd1 vccd1 vccd1 _06374_ sky130_fd_sc_hd__and3_1
X_14911_ net1317 vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_125_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12883__A1 _05756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15891_ net1364 vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_125_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11384__A team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17630_ clknet_leaf_3_wb_clk_i _03315_ _01571_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[16\]
+ sky130_fd_sc_hd__dfrtp_4
X_14842_ net1371 vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__inv_2
XANTENNA__14085__B1 _04265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17561_ clknet_leaf_89_wb_clk_i _03248_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_11985_ net1887 net296 net474 vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__mux2_1
X_14773_ net1276 vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10646__A0 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16512_ clknet_leaf_5_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[10\]
+ _00495_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13724_ net3187 _04108_ net2098 vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__a21oi_1
X_10936_ net555 _07069_ vssd1 vssd1 vccd1 vccd1 _07276_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17492_ clknet_leaf_67_wb_clk_i _03179_ _01475_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10110__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12927__B _03652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16443_ clknet_leaf_80_wb_clk_i _02197_ _00426_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12419__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10867_ _07205_ _07206_ vssd1 vssd1 vccd1 vccd1 _07207_ sky130_fd_sc_hd__or2_2
X_13655_ net988 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] _04087_ _04088_
+ vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12606_ net1948 net257 net397 vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__mux2_1
X_16374_ clknet_leaf_88_wb_clk_i _02128_ _00357_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[97\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13586_ _03912_ _04029_ _03903_ _03906_ vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__o211a_1
XANTENNA__09264__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10798_ net513 _05898_ _06779_ _06811_ net548 net537 vssd1 vssd1 vccd1 vccd1 _07138_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_27_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10949__A1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09803__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12537_ net2677 net265 net403 vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15325_ net1240 vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__inv_2
XANTENNA__09020__C net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12468_ net3023 net270 net413 vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__mux2_1
X_15256_ net1214 vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__inv_2
XANTENNA__09955__C net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11419_ _04478_ _07702_ vssd1 vssd1 vccd1 vccd1 _07733_ sky130_fd_sc_hd__nand2_1
X_14207_ net1753 vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12154__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15187_ net1419 vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__inv_2
X_12399_ net2125 net205 net419 vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__mux2_1
X_14138_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[127\] _04263_ _04267_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11993__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13115__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14069_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[92\] _04240_ _04249_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_33_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12874__A1 _05833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08630_ net376 vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__inv_2
X_17828_ clknet_leaf_91_wb_clk_i _03504_ _01768_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[98\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14076__B1 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08561_ net1077 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[19\] net940
+ vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__and3_1
X_17759_ clknet_leaf_98_wb_clk_i _03435_ _01699_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[29\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_81_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09699__A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08492_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[23\] net696 _04802_
+ _04805_ _04814_ vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_112_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_112_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_71_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12329__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09255__B1 _05593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08108__A _04504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09113_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[13\] net702 _05449_ _05452_
+ vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout316_A _07939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10076__C net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1058_A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09044_ net1107 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[12\] net937
+ vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__and3_1
XFILLER_0_142_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14000__B1 _04259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09558__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold420 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1955 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12064__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold431 team_01_WB.instance_to_wrap.a1.ADR_I\[20\] vssd1 vssd1 vccd1 vccd1 net1966
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10168__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold442 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1977 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1225_A net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold453 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1988 sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1999 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold475 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[8\] vssd1 vssd1 vccd1 vccd1
+ net2010 sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2021 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout900 net901 vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__buf_4
XANTENNA_fanout685_A _04780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold497 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2032 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout911 net913 vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__clkbuf_2
Xfanout922 _04770_ vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__buf_4
X_09946_ net998 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[3\] net959 vssd1
+ vssd1 vccd1 vccd1 _06286_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1013_X net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08778__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout933 _04765_ vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__buf_4
Xfanout944 _04756_ vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__buf_8
XANTENNA__13511__C1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout955 _04660_ vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_5_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout977 _04635_ vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__buf_6
Xhold1120 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[33\] vssd1 vssd1 vccd1 vccd1
+ net2655 sky130_fd_sc_hd__dlygate4sd3_1
X_09877_ _05416_ _06189_ vssd1 vssd1 vccd1 vccd1 _06217_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout852_A net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout473_X net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout988 net989 vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout999 net1003 vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08533__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1131 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2666 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1142 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2677 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08828_ net1105 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[1\] net894 vssd1
+ vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__and3_1
Xhold1153 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2688 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1164 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2699 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1175 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[104\] vssd1 vssd1 vccd1 vccd1
+ net2710 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1186 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2721 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1197 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2732 sky130_fd_sc_hd__dlygate4sd3_1
X_08759_ net1094 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[4\] net926 vssd1
+ vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout640_X net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout738_X net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10628__A0 _04706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ net2367 net270 net496 vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__mux2_1
XANTENNA__13290__A1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08944__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10721_ _07006_ _07013_ net534 vssd1 vssd1 vccd1 vccd1 _07061_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout905_X net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12239__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11143__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13440_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] _04945_ vssd1 vssd1
+ vccd1 vccd1 _03901_ sky130_fd_sc_hd__xnor2_1
X_10652_ net548 net513 vssd1 vssd1 vccd1 vccd1 _06992_ sky130_fd_sc_hd__or2_1
XANTENNA__09246__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13371_ _04517_ net565 net827 vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__o21a_1
X_10583_ _06901_ _06917_ vssd1 vssd1 vccd1 vccd1 _06923_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12322_ net2324 net315 net433 vssd1 vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15110_ net1381 vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_118_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16090_ clknet_leaf_132_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[12\]
+ _00078_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[12\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__08305__X _04645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15041_ net1280 vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__inv_2
X_12253_ net2169 net309 net440 vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11204_ _06218_ _07173_ _06194_ vssd1 vssd1 vccd1 vccd1 _07544_ sky130_fd_sc_hd__a21o_1
X_12184_ net2251 net294 net450 vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11135_ _07040_ _07338_ _07471_ net344 _07474_ vssd1 vssd1 vccd1 vccd1 _07475_ sky130_fd_sc_hd__o221a_1
XANTENNA__12702__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16992_ clknet_leaf_45_wb_clk_i _02679_ _00975_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11066_ _05491_ _06158_ _07366_ vssd1 vssd1 vccd1 vccd1 _07406_ sky130_fd_sc_hd__or3b_1
X_15943_ net1412 vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10017_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[1\] net757 _06355_ _06356_
+ vssd1 vssd1 vccd1 vccd1 _06357_ sky130_fd_sc_hd__a211o_1
X_15874_ net1229 vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__inv_2
XANTENNA__14058__B1 _04146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10331__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17613_ clknet_leaf_130_wb_clk_i _03298_ _01554_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14825_ net1294 vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09015__C net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17544_ clknet_leaf_63_wb_clk_i _03231_ _01527_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13281__A1 _07650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14756_ net1188 vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__inv_2
XANTENNA__09485__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11968_ net1793 net204 net471 vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__mux2_1
XANTENNA__08854__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13707_ net2375 _04100_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[2\]
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__12149__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10919_ _05374_ net339 vssd1 vssd1 vccd1 vccd1 _07259_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17475_ clknet_leaf_25_wb_clk_i _03162_ _01458_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_14687_ net1306 vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11899_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[25\] net207 net481 vssd1
+ vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__mux2_1
X_17945__1460 vssd1 vssd1 vccd1 vccd1 _17945__1460/HI net1460 sky130_fd_sc_hd__conb_1
XANTENNA__13569__C1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16426_ clknet_leaf_132_wb_clk_i _02180_ _00409_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13638_ net186 _04073_ _04074_ net725 vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__a211o_1
XANTENNA__09237__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11988__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16357_ clknet_leaf_122_wb_clk_i _02111_ _00340_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[80\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13569_ net185 _04015_ _04016_ net723 vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__a211o_1
XANTENNA__12792__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15308_ net1259 vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16288_ clknet_leaf_97_wb_clk_i _02042_ _00271_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11289__A team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15984__A net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15239_ net1390 vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_719 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09800_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[14\] net775 net735 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06140_ sky130_fd_sc_hd__a22o_1
XANTENNA__08763__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout207 net209 vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__buf_2
Xfanout218 _07831_ vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__buf_2
XANTENNA__12612__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout229 net232 vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__buf_2
X_07992_ net1097 vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09731_ net1132 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[20\] net975
+ vssd1 vssd1 vccd1 vccd1 _06071_ sky130_fd_sc_hd__and3_1
XANTENNA__10640__B _06928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10858__A0 _06158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09662_ _05999_ _06000_ vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__nand2_1
XANTENNA__14049__B1 _04258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08613_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[11\] net680 net667 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__a22o_1
X_09593_ _05707_ _05735_ vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__xnor2_2
X_08544_ _04883_ vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09476__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08475_ net1020 net880 vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__and2_1
XANTENNA__10368__A _06707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout433_A _07964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12059__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08109__Y _04579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1175_A team_01_WB.instance_to_wrap.cpu.DM0.dhit vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11898__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire619 _05315_ vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout600_A _04754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10389__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12783__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_80_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_32_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09027_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[9\] _04771_ _05344_ _05353_
+ _05355_ vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_131_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15894__A net1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1130_X net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12904__B1_N net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09892__A net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold250 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1785 sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1796 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09400__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout590_X net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout688_X net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold272 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1807 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 team_01_WB.instance_to_wrap.cpu.f0.write_data\[2\] vssd1 vssd1 vccd1 vccd1
+ net1818 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1829 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout730 net733 vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__clkbuf_8
Xfanout741 _04685_ vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08939__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09929_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[4\] net824 net790 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06269_ sky130_fd_sc_hd__a22o_1
Xfanout752 _04678_ vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08301__A net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout763 net764 vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__buf_2
Xfanout774 _04669_ vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__clkbuf_8
Xfanout785 net786 vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__clkbuf_8
Xfanout796 net797 vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__buf_4
XFILLER_0_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12940_ _05005_ _07757_ _03694_ vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__o21ai_1
X_12871_ net873 net378 vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__and2b_2
XFILLER_0_87_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14610_ net1308 vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__inv_2
X_11822_ net1958 net315 net493 vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15590_ net1383 vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__inv_2
XANTENNA__09467__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08674__C net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09132__A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11753_ net2845 net313 net500 vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__mux2_1
X_14541_ net1410 vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10704_ _05806_ net513 vssd1 vssd1 vccd1 vccd1 _07044_ sky130_fd_sc_hd__nor2_1
XANTENNA__09482__A3 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17260_ clknet_leaf_149_wb_clk_i _02947_ _01243_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14472_ net1347 vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__inv_2
X_11684_ net2166 net230 net501 vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16211_ clknet_leaf_124_wb_clk_i _01971_ _00199_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__dfrtp_1
XANTENNA__13566__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10635_ _04707_ _05835_ vssd1 vssd1 vccd1 vccd1 _06975_ sky130_fd_sc_hd__nor2_1
X_13423_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] net1170 net729 _04838_ net1127
+ vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__a32o_1
XFILLER_0_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17191_ clknet_leaf_104_wb_clk_i _02878_ _01174_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12774__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload109 clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload109/Y sky130_fd_sc_hd__clkinv_4
X_16142_ clknet_leaf_128_wb_clk_i _01905_ _00130_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13354_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[13\] _03826_ net827 vssd1 vssd1
+ vccd1 vccd1 _01881_ sky130_fd_sc_hd__mux2_1
X_10566_ net525 net521 vssd1 vssd1 vccd1 vccd1 _06906_ sky130_fd_sc_hd__nand2_4
XFILLER_0_140_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12305_ net2818 net233 net431 vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__mux2_1
X_13285_ _04621_ _03753_ _03772_ net825 vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__o31a_1
X_16073_ clknet_leaf_152_wb_clk_i _01866_ _00061_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\]
+ sky130_fd_sc_hd__dfstp_2
X_10497_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[31\] net799 net782 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06837_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10444__C net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15024_ net1276 vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__inv_2
X_12236_ net2979 net241 net441 vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__mux2_1
XANTENNA__12432__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12167_ net1845 net200 net448 vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__mux2_1
X_11118_ _06928_ _07133_ _07457_ net328 vssd1 vssd1 vccd1 vccd1 _07458_ sky130_fd_sc_hd__a211o_1
XANTENNA__12829__A1 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12098_ net2615 net206 net457 vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__mux2_1
X_16975_ clknet_leaf_33_wb_clk_i _02662_ _00958_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_15926_ net1415 vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__inv_2
X_11049_ net517 _06339_ vssd1 vssd1 vccd1 vccd1 _07389_ sky130_fd_sc_hd__or2_1
Xinput7 DAT_I[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10304__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15857_ net1344 vssd1 vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__inv_2
XFILLER_0_149_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14808_ net1215 vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09458__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15788_ net1190 vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08584__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17527_ clknet_leaf_13_wb_clk_i _03214_ _01510_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_14739_ net1194 vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__inv_2
XANTENNA__14883__A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08260_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[21\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[13\]
+ net1050 vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__mux2_1
X_17458_ clknet_leaf_145_wb_clk_i _03145_ _01441_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08881__A net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16409_ clknet_leaf_124_wb_clk_i _02163_ _00392_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_08191_ net2838 net2448 net1052 vssd1 vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12607__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17389_ clknet_leaf_109_wb_clk_i _03076_ _01372_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12765__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11511__S net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10635__B _05835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08984__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_93_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13190__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08736__A2 _05074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12342__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08759__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07975_ team_01_WB.instance_to_wrap.cpu.f0.i\[21\] vssd1 vssd1 vccd1 vccd1 _04473_
+ sky130_fd_sc_hd__inv_2
XANTENNA__10370__B _05566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout383_A _03570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16111__Q team_01_WB.instance_to_wrap.cpu.f0.data_adr\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09714_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[21\] net812 net773 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[21\]
+ _06053_ vssd1 vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__a221o_1
X_09645_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[23\] net817 net791 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[23\]
+ _05984_ vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout550_A _05151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1292_A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout648_A _04823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09576_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[25\] net802 _05904_
+ _05911_ _05913_ vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_78_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09449__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13245__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_33_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08527_ net1001 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[18\] net910
+ vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1080_X net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout815_A net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout436_X net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1178_X net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09887__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08458_ net1081 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[23\] net891
+ vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08791__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13548__A2 _07154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12517__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08389_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[2\] _04623_ _04626_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_34_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout603_X net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12756__B1 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10420_ net1132 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[27\] net945
+ vssd1 vssd1 vccd1 vccd1 _06760_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_154_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08975__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10351_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[17\] net819 net744 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _06691_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_111_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13070_ net2750 net2647 net852 vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__mux2_1
XANTENNA__13856__B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10282_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[19\] net817 net772 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _06622_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout972_X net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12021_ net2196 net305 net469 vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08727__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15129__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10561__A _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12252__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10534__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08669__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout560 net561 vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11166__A1_N net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout571 net572 vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__clkbuf_2
XANTENNA__14130__C1 net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16760_ clknet_leaf_61_wb_clk_i _02447_ _00743_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout593 _04845_ vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__clkbuf_4
X_13972_ _04222_ _04237_ _04239_ vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__and3_4
XANTENNA__08966__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10298__A1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15711_ net1317 vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__inv_2
X_12923_ net1579 net869 net356 _03691_ vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__a22o_1
X_16691_ clknet_leaf_20_wb_clk_i _02378_ _00674_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_15642_ net1373 vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__inv_2
X_12854_ net2167 net225 net379 vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11805_ net3115 net233 net491 vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15573_ net1276 vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12785_ net1725 net638 net606 _03618_ vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17312_ clknet_leaf_47_wb_clk_i _02999_ _01295_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09797__A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14524_ net1407 vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_1_Left_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11736_ net1898 net293 net500 vssd1 vssd1 vccd1 vccd1 _03220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12935__B net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17243_ clknet_leaf_70_wb_clk_i _02930_ _01226_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14455_ net1227 vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__inv_2
X_11667_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[18\] _07251_ net713 vssd1 vssd1
+ vccd1 vccd1 _07871_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12427__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12747__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13406_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\] net596 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10618_ _06950_ _06957_ net520 vssd1 vssd1 vccd1 vccd1 _06958_ sky130_fd_sc_hd__mux2_1
X_17174_ clknet_leaf_30_wb_clk_i _02861_ _01157_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14386_ net1193 vssd1 vssd1 vccd1 vccd1 _00180_ sky130_fd_sc_hd__inv_2
X_11598_ _07814_ vssd1 vssd1 vccd1 vccd1 _07815_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_12_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire961 _04656_ vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10222__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16125_ clknet_leaf_124_wb_clk_i _00025_ _00113_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__dfrtp_1
Xwire983 _04631_ vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10549_ net510 net509 net543 vssd1 vssd1 vccd1 vccd1 _06889_ sky130_fd_sc_hd__mux2_1
X_13337_ net1071 _07682_ _03811_ _04518_ vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__a211o_1
XFILLER_0_51_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16056_ clknet_leaf_150_wb_clk_i _01849_ _00044_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_13268_ team_01_WB.instance_to_wrap.cpu.f0.i\[28\] _03749_ vssd1 vssd1 vccd1 vccd1
+ _03759_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15007_ net1318 vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__inv_2
X_12219_ net2420 net308 net446 vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__mux2_1
XANTENNA__12162__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13199_ net9 net836 net628 net1655 vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__o22a_1
XANTENNA__11722__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11286__B _07056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16958_ clknet_leaf_85_wb_clk_i _02645_ _00941_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09143__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15909_ net1417 vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__inv_2
X_16889_ clknet_leaf_104_wb_clk_i _02576_ _00872_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09430_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[28\] net700 net654 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13227__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_149_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09361_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[25\] net671 net668 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[25\]
+ _05685_ vssd1 vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__a221o_1
XANTENNA__09203__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08312_ net1137 net984 vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__and2_1
XANTENNA__10349__C net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_19_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09292_ net1084 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[22\] net918
+ vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17697__Q team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_75_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_12 _03663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_7_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08243_ net2585 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[30\] net1042 vssd1 vssd1
+ vccd1 vccd1 _03444_ sky130_fd_sc_hd__mux2_1
XANTENNA__09500__A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_34 net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12337__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12738__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09879__A_N net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_45 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_56 _03654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout229_A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08174_ net1748 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[99\] net1054 vssd1 vssd1
+ vccd1 vccd1 _03513_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_132_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08116__A team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_144_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16106__Q team_01_WB.instance_to_wrap.cpu.f0.data_adr\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08957__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1040_A net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10764__A2 _06811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1138_A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput130 net130 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__buf_2
Xoutput141 net141 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__buf_2
XANTENNA_fanout598_A net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13163__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput152 net152 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
Xoutput163 net163 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__clkbuf_4
Xoutput174 net174 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__clkbuf_4
X_18018__1512 vssd1 vssd1 vccd1 vccd1 _18018__1512/HI net1512 sky130_fd_sc_hd__conb_1
XANTENNA__12072__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11713__A1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10516__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09382__A2 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout386_X net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout765_A net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08590__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08786__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout932_A net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09628_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[23\] net794 net739 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_52_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout720_X net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09559_ _05898_ vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout818_X net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12570_ net2120 net267 net400 vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09842__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12755__B team_01_WB.instance_to_wrap.cpu.f0.data_adr\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11521_ net1173 _07784_ vssd1 vssd1 vccd1 vccd1 _07785_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12247__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14240_ net1189 vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__inv_2
X_11452_ _07672_ _07750_ vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10403_ _06641_ _06677_ _06715_ _06742_ vssd1 vssd1 vccd1 vccd1 _06743_ sky130_fd_sc_hd__or4_1
X_14171_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[7\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[6\]
+ _04189_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__and3_1
XANTENNA__11401__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11383_ team_01_WB.instance_to_wrap.cpu.f0.i\[22\] _07700_ _07710_ vssd1 vssd1 vccd1
+ vccd1 _07712_ sky130_fd_sc_hd__and3_1
XANTENNA__11952__A1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10334_ net559 _05568_ _04883_ vssd1 vssd1 vccd1 vccd1 _06674_ sky130_fd_sc_hd__o21ai_1
XANTENNA_input61_A wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13122_ net1604 net843 net632 team_01_WB.instance_to_wrap.a1.ADR_I\[21\] vssd1 vssd1
+ vccd1 vccd1 _02019_ sky130_fd_sc_hd__a22o_1
XANTENNA__08313__X _04653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13154__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17930_ net1447 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
X_13053_ net2655 net2553 net865 vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__mux2_1
XANTENNA__10291__A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10265_ net1128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[19\] net945
+ vssd1 vssd1 vccd1 vccd1 _06605_ sky130_fd_sc_hd__and3_1
Xfanout1300 net1301 vssd1 vssd1 vccd1 vccd1 net1300 sky130_fd_sc_hd__buf_2
XANTENNA__12901__B1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12004_ net2819 net270 net468 vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__mux2_1
Xfanout1311 net1322 vssd1 vssd1 vccd1 vccd1 net1311 sky130_fd_sc_hd__buf_4
X_17861_ clknet_leaf_126_wb_clk_i _03536_ _01801_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09373__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10196_ net992 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[8\] net954 vssd1
+ vssd1 vccd1 vccd1 _06536_ sky130_fd_sc_hd__and3_1
Xfanout1322 net1430 vssd1 vssd1 vccd1 vccd1 net1322 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_139_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1333 net1334 vssd1 vssd1 vccd1 vccd1 net1333 sky130_fd_sc_hd__buf_4
XANTENNA__11674__X _07877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1344 net1430 vssd1 vssd1 vccd1 vccd1 net1344 sky130_fd_sc_hd__buf_2
XFILLER_0_108_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16812_ clknet_leaf_147_wb_clk_i _02499_ _00795_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1355 net1369 vssd1 vssd1 vccd1 vccd1 net1355 sky130_fd_sc_hd__buf_2
Xfanout1366 net1368 vssd1 vssd1 vccd1 vccd1 net1366 sky130_fd_sc_hd__buf_4
XANTENNA__12710__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17792_ clknet_leaf_117_wb_clk_i net2726 _01732_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_128_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_91_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1377 net1429 vssd1 vssd1 vccd1 vccd1 net1377 sky130_fd_sc_hd__buf_2
Xfanout1388 net1391 vssd1 vssd1 vccd1 vccd1 net1388 sky130_fd_sc_hd__buf_4
Xfanout390 _03569_ vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_128_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1399 net1409 vssd1 vssd1 vccd1 vccd1 net1399 sky130_fd_sc_hd__buf_4
XFILLER_0_89_915 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11468__B1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16743_ clknet_leaf_106_wb_clk_i _02430_ _00726_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13955_ _04219_ _04222_ _04237_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__and3_4
X_12906_ net1904 net872 net359 _03679_ vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__a22o_1
XANTENNA__13107__A net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16674_ clknet_leaf_76_wb_clk_i _02361_ _00657_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13886_ _04190_ _04191_ _04192_ vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__or3_1
XANTENNA__10140__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08884__B2 net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15625_ net1296 vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12837_ net2646 net214 net380 vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15556_ net1230 vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__inv_2
XANTENNA__09833__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12768_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] net1061 net362 _03606_
+ vssd1 vssd1 vccd1 vccd1 _03607_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08862__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14507_ net1415 vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11719_ net1819 net300 net499 vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__mux2_1
X_15487_ net1318 vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12699_ net2123 net271 net385 vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17226_ clknet_leaf_11_wb_clk_i _02913_ _01209_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14438_ net1307 vssd1 vssd1 vccd1 vccd1 _00232_ sky130_fd_sc_hd__inv_2
Xinput10 DAT_I[17] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
Xinput21 DAT_I[27] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput32 DAT_I[8] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
Xinput43 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11996__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput54 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_1
X_17157_ clknet_leaf_51_wb_clk_i _02844_ _01140_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold805 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2340 sky130_fd_sc_hd__dlygate4sd3_1
Xinput65 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_1
X_14369_ net1208 vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold816 _03520_ vssd1 vssd1 vccd1 vccd1 net2351 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold827 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2362 sky130_fd_sc_hd__dlygate4sd3_1
X_16108_ clknet_leaf_137_wb_clk_i _01883_ _00096_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[15\]
+ sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_137_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_137_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold838 _03456_ vssd1 vssd1 vccd1 vccd1 net2373 sky130_fd_sc_hd__dlygate4sd3_1
X_17088_ clknet_leaf_48_wb_clk_i _02775_ _01071_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold849 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2384 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13145__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08930_ net1028 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[6\] net924 vssd1
+ vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__and3_1
X_16039_ clknet_leaf_88_wb_clk_i _01833_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08861_ net1017 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[3\] net927 vssd1
+ vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_36_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1505 team_01_WB.instance_to_wrap.cpu.f0.num\[26\] vssd1 vssd1 vccd1 vccd1 net3040
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1516 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[15\] vssd1 vssd1 vccd1 vccd1
+ net3051 sky130_fd_sc_hd__dlygate4sd3_1
X_08792_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[0\] net671 _05129_ _05130_
+ _05131_ vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12620__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1527 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net3062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1538 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1 net3073
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_88_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1549 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[11\] vssd1 vssd1 vccd1 vccd1
+ net3084 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_88_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09413_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[27\] net676 net652 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[27\]
+ _05739_ vssd1 vssd1 vccd1 vccd1 _05753_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10079__C net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout346_A net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1088_A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09344_ net1115 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[25\] net909
+ vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_62_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09230__A net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09275_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[20\] net701 _05610_ _05614_
+ vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__o22a_2
XFILLER_0_75_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10376__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12067__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_136_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1255_A net1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08226_ net2828 net2774 net1048 vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_151_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13958__Y _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16501__CLK clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08157_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[124\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[116\]
+ net1045 vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08088_ _04525_ _04559_ _04560_ net569 net1578 vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout882_A net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13136__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13974__X _04266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10050_ _06386_ _06387_ _06388_ _06389_ vssd1 vssd1 vccd1 vccd1 _06390_ sky130_fd_sc_hd__or4_1
XANTENNA__09355__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout670_X net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout768_X net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12530__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08947__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09107__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14100__A2 _04226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout935_X net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_82_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13740_ net1178 net1065 net1539 vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__a21o_1
XANTENNA__10122__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10952_ _06255_ _06410_ _07291_ _06468_ vssd1 vssd1 vccd1 vccd1 _07292_ sky130_fd_sc_hd__a31o_1
XFILLER_0_86_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_123_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13671_ net1625 net568 net347 team_01_WB.instance_to_wrap.cpu.f0.i\[30\] vssd1 vssd1
+ vccd1 vccd1 _01831_ sky130_fd_sc_hd__a22o_1
X_10883_ _05566_ _06707_ vssd1 vssd1 vccd1 vccd1 _07223_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08963__B net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15410_ net1291 vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12622_ net2977 net188 net391 vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__mux2_1
X_16390_ clknet_leaf_88_wb_clk_i net2643 _00373_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[113\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09815__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08308__X _04648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08682__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15341_ net1266 vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12553_ net2114 net315 net404 vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11504_ net1726 net876 _07758_ _07779_ vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__o22a_1
XFILLER_0_124_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15272_ net1387 vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12484_ net1999 net312 net414 vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_91_Left_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17011_ clknet_leaf_16_wb_clk_i _02698_ _00994_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_14223_ net3127 vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11669__X _07873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11435_ team_01_WB.instance_to_wrap.cpu.f0.i\[9\] _07736_ net324 vssd1 vssd1 vccd1
+ vccd1 _07742_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12705__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input64_X net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11366_ team_01_WB.instance_to_wrap.cpu.f0.i\[24\] team_01_WB.instance_to_wrap.cpu.f0.i\[23\]
+ net1069 _07694_ vssd1 vssd1 vccd1 vccd1 _07695_ sky130_fd_sc_hd__and4_1
X_14154_ net1583 net605 _04437_ net1183 vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10733__B _05898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13105_ _03723_ _03724_ _03725_ _03728_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__or4_4
X_10317_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[18\] net730 _06654_ _06655_
+ _06656_ vssd1 vssd1 vccd1 vccd1 _06657_ sky130_fd_sc_hd__a2111o_1
X_11297_ net199 net195 _07635_ vssd1 vssd1 vccd1 vccd1 _07637_ sky130_fd_sc_hd__o21ai_1
X_14085_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[100\] _04254_ _04265_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[4\]
+ _04372_ vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__a221o_1
XANTENNA__10452__C net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09346__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17913_ net1444 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
X_10248_ net768 _06572_ _06575_ _06587_ vssd1 vssd1 vccd1 vccd1 _06588_ sky130_fd_sc_hd__or4_1
X_13036_ net2222 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[58\] net863 vssd1 vssd1
+ vccd1 vccd1 _02089_ sky130_fd_sc_hd__mux2_1
XANTENNA__09018__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1130 net1134 vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__clkbuf_2
Xfanout1141 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[19\] vssd1 vssd1 vccd1 vccd1
+ net1141 sky130_fd_sc_hd__buf_2
X_17844_ clknet_leaf_91_wb_clk_i net2351 _01784_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[114\]
+ sky130_fd_sc_hd__dfrtp_1
X_10179_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[10\] net796 net761 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[10\]
+ _06518_ vssd1 vssd1 vccd1 vccd1 _06519_ sky130_fd_sc_hd__a221o_1
XANTENNA__12440__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1152 net1153 vssd1 vssd1 vccd1 vccd1 net1152 sky130_fd_sc_hd__buf_2
Xfanout1163 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[17\] vssd1 vssd1 vccd1 vccd1
+ net1163 sky130_fd_sc_hd__buf_2
Xfanout1174 team_01_WB.instance_to_wrap.cpu.DM0.ihit vssd1 vssd1 vccd1 vccd1 net1174
+ sky130_fd_sc_hd__buf_2
Xfanout1185 _00026_ vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08857__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1196 net1201 vssd1 vssd1 vccd1 vccd1 net1196 sky130_fd_sc_hd__buf_2
X_17775_ clknet_leaf_101_wb_clk_i _03451_ _01715_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[45\]
+ sky130_fd_sc_hd__dfstp_1
X_14987_ net1423 vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__inv_2
X_16726_ clknet_leaf_29_wb_clk_i _02413_ _00709_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11283__C _07553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13938_ _04225_ _04229_ vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__nor2_4
XFILLER_0_44_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16657_ clknet_leaf_116_wb_clk_i _02344_ _00640_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10748__X _07088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13869_ net1177 net1064 net2427 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[30\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_29_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18009__1509 vssd1 vssd1 vccd1 vccd1 _18009__1509/HI net1509 sky130_fd_sc_hd__conb_1
X_15608_ net1209 vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__inv_2
XFILLER_0_147_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09806__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13602__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16588_ clknet_leaf_148_wb_clk_i _02275_ _00571_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15539_ net1392 vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__inv_2
XANTENNA__11613__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14891__A net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09060_ net1029 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[12\] net907
+ vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12169__A1 _07866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08011_ team_01_WB.instance_to_wrap.a1.READ_I vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__inv_2
XANTENNA__13366__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17209_ clknet_leaf_100_wb_clk_i _02896_ _01192_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09034__A1 _05373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12615__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold602 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold613 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2148 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13300__A net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold624 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2159 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold635 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2170 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold646 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2181 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13118__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold657 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2203 sky130_fd_sc_hd__dlygate4sd3_1
X_09962_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[3\] net800 net792 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06302_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold679 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2214 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08913_ _05249_ _05250_ _05251_ _05252_ vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_139_Left_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09893_ net1152 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[5\] net955 vssd1
+ vssd1 vccd1 vccd1 _06233_ sky130_fd_sc_hd__and3_1
XFILLER_0_85_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1302 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2837 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12350__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1313 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2848 sky130_fd_sc_hd__dlygate4sd3_1
X_08844_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[1\] net652 _05165_ _05169_
+ _05172_ vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10352__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1324 _02141_ vssd1 vssd1 vccd1 vccd1 net2859 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1003_A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1335 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1346 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2881 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1357 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2892 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1368 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[12\] vssd1 vssd1 vccd1 vccd1
+ net2903 sky130_fd_sc_hd__dlygate4sd3_1
X_08775_ net598 _05110_ _05113_ vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout463_A _07954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1379 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2914 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_34_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_0_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10655__A1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout630_A _03738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09598__C net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09327_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[24\] net665 _04808_
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[24\] _05666_ vssd1 vssd1 vccd1
+ vccd1 _05667_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1160_X net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout516_X net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1258_X net1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10958__A2 _06924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14149__A2 _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09258_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[20\] net699 net670 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08209_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[72\] net2945 net1046 vssd1 vssd1
+ vccd1 vccd1 _03478_ sky130_fd_sc_hd__mux2_1
X_09189_ _05495_ _05528_ net600 vssd1 vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__mux2_2
XANTENNA__12525__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11220_ net368 _07343_ _07344_ net335 _07559_ vssd1 vssd1 vccd1 vccd1 _07560_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_79_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09576__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08304__A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout885_X net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11151_ _07449_ net321 _07490_ vssd1 vssd1 vccd1 vccd1 _07491_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10102_ _06441_ vssd1 vssd1 vccd1 vccd1 _06442_ sky130_fd_sc_hd__inv_2
XANTENNA__09328__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11082_ _04844_ _05997_ _07418_ _07419_ _07421_ vssd1 vssd1 vccd1 vccd1 _07422_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12868__C1 _03652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10033_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[0\] net815 net734 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06373_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_8_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14910_ net1345 vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__inv_2
XANTENNA__12260__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15890_ net1347 vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__inv_2
XANTENNA__12883__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08677__C net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input24_A DAT_I[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14841_ net1231 vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17560_ clknet_leaf_89_wb_clk_i _03247_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_19_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14772_ net1378 vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__inv_2
X_11984_ net1940 net279 net472 vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__mux2_1
XANTENNA__08974__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16511_ clknet_leaf_5_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[9\]
+ _00494_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10646__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13723_ net2423 _04108_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[13\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_105_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10935_ net558 _07069_ vssd1 vssd1 vccd1 vccd1 _07275_ sky130_fd_sc_hd__and2_1
X_17491_ clknet_leaf_18_wb_clk_i _03178_ _01474_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16442_ clknet_leaf_69_wb_clk_i _02196_ _00425_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13654_ net727 _07449_ net988 vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_155_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10866_ net562 _07192_ _07193_ _07203_ net555 vssd1 vssd1 vccd1 vccd1 _07206_ sky130_fd_sc_hd__a32o_1
XFILLER_0_85_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12605_ net2334 net229 net397 vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__mux2_1
X_16373_ clknet_leaf_122_wb_clk_i _02127_ _00356_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[96\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09301__C net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13585_ _03912_ _04029_ _03906_ vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__o21ai_1
X_10797_ _05931_ _05963_ net510 net509 net549 net536 vssd1 vssd1 vccd1 vccd1 _07137_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10447__C _04660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15324_ net1245 vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__inv_2
XFILLER_0_147_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12536_ net3018 net233 net403 vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15255_ net1244 vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12435__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12467_ net2476 net242 net413 vssd1 vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_144_Right_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14206_ net2257 vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__clkbuf_1
X_11418_ _07691_ _07732_ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__nor2_1
X_15186_ net1292 vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12398_ net2434 net272 net421 vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14137_ _04416_ _04417_ _04419_ _04421_ vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__or4_1
X_11349_ team_01_WB.instance_to_wrap.cpu.f0.i\[11\] _07677_ vssd1 vssd1 vccd1 vccd1
+ _07678_ sky130_fd_sc_hd__nand2_2
XANTENNA__08501__X _04841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14068_ net3125 net604 vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__or2_1
X_17908__1519 vssd1 vssd1 vccd1 vccd1 net1519 _17908__1519/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_33_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13870__A_N net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12170__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13019_ net2490 net2336 net861 vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__mux2_1
XANTENNA__12874__A2 _07752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10885__A1 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08587__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17827_ clknet_leaf_93_wb_clk_i _03503_ _01767_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[97\]
+ sky130_fd_sc_hd__dfrtp_1
X_08560_ _04889_ _04893_ _04895_ _04899_ vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__or4_1
X_17758_ clknet_leaf_99_wb_clk_i _03434_ _01698_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[28\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10637__A1 _05835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16709_ clknet_leaf_51_wb_clk_i _02396_ _00692_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_08491_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[23\] net670 _04812_ _04820_
+ _04798_ vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__a2111o_1
X_17689_ clknet_leaf_128_wb_clk_i _03373_ _01630_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_49_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11514__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09211__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09255__A1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08058__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09112_ _05443_ _05444_ _05450_ _05451_ vssd1 vssd1 vccd1 vccd1 _05452_ sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_152_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_152_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_143_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13339__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10925__Y _07265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09043_ net1111 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[12\] net908
+ vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14000__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12345__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout211_A net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold410 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1945 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09558__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold421 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net1956 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold432 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1967 sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1978 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16114__Q team_01_WB.instance_to_wrap.cpu.f0.data_adr\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold454 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net1989 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_147_Left_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1120_A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold465 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2000 sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 _03339_ vssd1 vssd1 vccd1 vccd1 net2011 sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2022 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout901 _04788_ vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_74_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold498 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2033 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout912 net913 vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__buf_4
X_09945_ _06280_ _06283_ vssd1 vssd1 vccd1 vccd1 _06285_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout923 _04770_ vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout580_A _07752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12314__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout934 net935 vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_146_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout678_A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout945 net946 vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12080__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09226__Y _05566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout956 net957 vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] _06215_ net623 vssd1
+ vssd1 vccd1 vccd1 _06216_ sky130_fd_sc_hd__mux2_2
Xhold1110 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2645 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout989 _04499_ vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__buf_4
Xhold1121 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2656 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1132 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2667 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08827_ net1106 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[1\] net903 vssd1
+ vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__and3_1
XANTENNA__13971__Y _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1143 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[71\] vssd1 vssd1 vccd1 vccd1
+ net2678 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14796__A net1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout466_X net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout845_A net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1154 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2689 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1165 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2700 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1176 _02143_ vssd1 vssd1 vccd1 vccd1 net2711 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1187 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2722 sky130_fd_sc_hd__dlygate4sd3_1
X_08758_ net1099 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[4\] net912 vssd1
+ vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__and3_1
XANTENNA__08794__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1198 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2733 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_120_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10628__A1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_156_Left_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08689_ net1008 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[7\] net934 vssd1
+ vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__and3_1
XANTENNA__09494__A1 team_01_WB.instance_to_wrap.cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout633_X net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10720_ _07058_ _07059_ net517 vssd1 vssd1 vccd1 vccd1 _07060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09121__C net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout800_X net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10651_ _06989_ _06990_ net536 vssd1 vssd1 vccd1 vccd1 _06991_ sky130_fd_sc_hd__mux2_1
XANTENNA__10267__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10582_ net503 _06920_ vssd1 vssd1 vccd1 vccd1 _06922_ sky130_fd_sc_hd__nand2_1
X_13370_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[8\] net827 _07650_ _03837_ vssd1
+ vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__o22a_1
XFILLER_0_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12321_ net2611 net319 net434 vssd1 vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_118_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12255__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15040_ net1233 vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__inv_2
XANTENNA__09549__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12252_ net2902 net292 net441 vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__mux2_1
X_11203_ _06194_ _06218_ _07173_ vssd1 vssd1 vccd1 vccd1 _07543_ sky130_fd_sc_hd__nand3_1
X_12183_ net2785 net296 net450 vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08969__A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11134_ _07472_ _07473_ _07432_ vssd1 vssd1 vccd1 vccd1 _07474_ sky130_fd_sc_hd__a21o_1
X_16991_ clknet_leaf_39_wb_clk_i _02678_ _00974_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13502__B1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11395__A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15942_ net1407 vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__inv_2
X_11065_ _05454_ net373 _07371_ _07404_ vssd1 vssd1 vccd1 vccd1 _07405_ sky130_fd_sc_hd__a2bb2o_1
X_10016_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[1\] net737 net735 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06356_ sky130_fd_sc_hd__a22o_1
XANTENNA__09721__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15873_ net1229 vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__inv_2
XANTENNA_output130_A net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14824_ net1375 vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__inv_2
X_17612_ clknet_leaf_130_wb_clk_i _03297_ _01553_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10619__A1 _06958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17543_ clknet_leaf_107_wb_clk_i _03230_ _01526_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_14755_ net1202 vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__inv_2
X_11967_ net2584 net272 net473 vssd1 vssd1 vccd1 vccd1 _03015_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13706_ _04101_ _04123_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[3\]
+ sky130_fd_sc_hd__and2b_1
XANTENNA__11292__A1 net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17474_ clknet_leaf_76_wb_clk_i _03161_ _01457_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10918_ _04738_ _06591_ _06917_ _05374_ _04736_ vssd1 vssd1 vccd1 vccd1 _07258_ sky130_fd_sc_hd__a2111oi_1
X_14686_ net1227 vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11898_ net2185 net248 net481 vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16425_ clknet_leaf_140_wb_clk_i _02179_ _00408_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13637_ net197 net193 _07916_ net643 vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__o211a_1
X_10849_ _06469_ _06472_ _06568_ vssd1 vssd1 vccd1 vccd1 _07189_ sky130_fd_sc_hd__or3_1
XFILLER_0_156_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16356_ clknet_leaf_97_wb_clk_i net2679 _00339_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[79\]
+ sky130_fd_sc_hd__dfrtp_1
X_13568_ net196 net192 _07872_ net642 vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15307_ net1395 vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12792__A1 _07520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12519_ net2478 net317 net410 vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__mux2_1
X_16287_ clknet_leaf_92_wb_clk_i _02041_ _00270_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10474__A _06811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12165__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13499_ _03841_ _03951_ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_140_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15238_ net1404 vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_2_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13741__B1 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15169_ net1280 vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout208 net209 vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09960__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout219 net220 vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__buf_2
X_07991_ team_01_WB.instance_to_wrap.cpu.f0.i\[0\] vssd1 vssd1 vccd1 vccd1 _04489_
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_52_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09730_ net1145 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[20\] net979
+ vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__and3_1
XANTENNA__10858__A1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09661_ _05999_ _06000_ vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__and2_1
XANTENNA__09206__C net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08612_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[11\] net650 net648 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[11\]
+ _04951_ vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__a221o_1
X_09592_ net512 vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09503__A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08543_ net597 _04881_ _04882_ vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_82_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09997__X _06337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08474_ net1083 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[23\] net910
+ vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16109__Q team_01_WB.instance_to_wrap.cpu.f0.data_adr\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09779__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13980__B1 _04259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12075__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09026_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[9\] net680 _05343_ _05349_
+ _05360_ vssd1 vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_27_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13966__Y _04258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout795_A net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold240 _02029_ vssd1 vssd1 vccd1 vccd1 net1775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1786 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 team_01_WB.instance_to_wrap.a1.ADR_I\[28\] vssd1 vssd1 vccd1 vccd1 net1797
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_72_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold273 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1808 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10010__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold284 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1819 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold295 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1830 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout720 net722 vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__clkbuf_4
Xfanout731 net733 vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__clkbuf_8
X_09928_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[4\] net819 net784 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06268_ sky130_fd_sc_hd__a22o_1
Xfanout742 net744 vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__clkbuf_8
Xfanout753 net754 vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13496__C1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout764 net767 vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08301__B net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout775 _04667_ vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_137_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout786 _04659_ vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__buf_6
Xfanout797 _04651_ vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__buf_4
XANTENNA_fanout750_X net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09859_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[12\] net818 _04678_
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[12\] vssd1 vssd1 vccd1 vccd1
+ _06199_ sky130_fd_sc_hd__a22o_1
XANTENNA__11510__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15415__A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12870_ _04510_ _03575_ _03578_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_write_i
+ sky130_fd_sc_hd__nor3b_1
XFILLER_0_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11821_ net2804 net318 net494 vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14540_ net1421 vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__inv_2
X_11752_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] _07938_ net615 vssd1
+ vssd1 vccd1 vccd1 _07939_ sky130_fd_sc_hd__mux2_2
XFILLER_0_56_718 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10703_ _07038_ _07042_ net529 vssd1 vssd1 vccd1 vccd1 _07043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14471_ net1347 vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__inv_2
X_11683_ net612 _07811_ _07883_ _07882_ vssd1 vssd1 vccd1 vccd1 _07884_ sky130_fd_sc_hd__a31o_2
XANTENNA__08690__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16210_ clknet_leaf_123_wb_clk_i net1657 _00198_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__dfrtp_1
X_17907__1518 vssd1 vssd1 vccd1 vccd1 net1518 _17907__1518/LO sky130_fd_sc_hd__conb_1
X_13422_ _03861_ _03882_ _03860_ vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__a21oi_1
X_17190_ clknet_leaf_72_wb_clk_i _02877_ _01173_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10634_ _04707_ _05835_ vssd1 vssd1 vccd1 vccd1 _06974_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16141_ clknet_leaf_129_wb_clk_i _01904_ _00129_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13353_ net565 _07678_ _03823_ _03825_ net586 vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__a32o_1
X_10565_ net531 net516 vssd1 vssd1 vccd1 vccd1 _06905_ sky130_fd_sc_hd__nor2_2
XFILLER_0_107_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10785__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12304_ net2442 net239 net431 vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__mux2_1
X_16072_ clknet_leaf_152_wb_clk_i _01865_ _00060_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_122_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13284_ _04470_ _03752_ vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__and2_1
X_10496_ net1131 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[31\] net945
+ vssd1 vssd1 vccd1 vccd1 _06836_ sky130_fd_sc_hd__and3_1
X_15023_ net1388 vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12235_ net1942 net201 net439 vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__mux2_1
XANTENNA__12713__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10537__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12166_ net2605 net205 net447 vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__mux2_1
X_11117_ _06921_ _07121_ vssd1 vssd1 vccd1 vccd1 _07457_ sky130_fd_sc_hd__nor2_1
X_16974_ clknet_leaf_37_wb_clk_i _02661_ _00957_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12829__A2 _07476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12097_ net2450 net248 net457 vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__mux2_1
X_15925_ net1417 vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__inv_2
X_11048_ _07386_ _07387_ vssd1 vssd1 vccd1 vccd1 _07388_ sky130_fd_sc_hd__and2_1
Xinput8 DAT_I[15] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08363__D1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15856_ net1334 vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08865__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14807_ net1243 vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15787_ net1190 vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__inv_2
X_12999_ net2568 net2477 net856 vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14738_ net1194 vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__inv_2
X_17526_ clknet_leaf_30_wb_clk_i _03213_ _01509_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11999__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17457_ clknet_leaf_117_wb_clk_i _03144_ _01440_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_14669_ net1226 vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08881__B _05220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16408_ clknet_leaf_125_wb_clk_i _02162_ _00391_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_08190_ net2236 net2407 net1054 vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__mux2_1
X_17388_ clknet_leaf_146_wb_clk_i _03075_ _01371_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12765__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16339_ clknet_leaf_117_wb_clk_i net2630 _00322_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10240__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18009_ net1509 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__buf_2
XANTENNA__12623__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10932__A _05338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10528__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09933__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08402__A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07974_ team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1 vccd1 vccd1 _04472_
+ sky130_fd_sc_hd__inv_2
X_09713_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[21\] net785 net751 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__a22o_1
X_09644_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[23\] net821 net759 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05984_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09575_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[25\] net746 net740 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout543_A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_42_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1285_A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08526_ net1000 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[18\] net887 vssd1
+ vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__and3_1
XANTENNA__11256__B2 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08457_ net1112 net894 vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__and2_4
XFILLER_0_136_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout331_X net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout710_A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout808_A net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1073_X net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout429_X net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08388_ net1170 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[4\] _04624_ vssd1 vssd1
+ vccd1 vccd1 _04728_ sky130_fd_sc_hd__and3b_1
XANTENNA__12756__A1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12756__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10231__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10350_ net1139 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[17\] net955
+ vssd1 vssd1 vccd1 vccd1 _06690_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout798_X net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09009_ net1013 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[9\] net930 vssd1
+ vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__and3_1
XFILLER_0_143_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10281_ _06608_ _06612_ _06616_ _06620_ vssd1 vssd1 vccd1 vccd1 _06621_ sky130_fd_sc_hd__or4_1
XFILLER_0_104_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10519__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12533__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12020_ net2706 net310 net469 vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__mux2_1
XANTENNA__11657__B net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08312__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10561__B _04738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout965_X net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout550 _05151_ vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_81_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout561 _04749_ vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__clkbuf_4
Xfanout572 _04196_ vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13872__B net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13971_ _04218_ _04248_ vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__nor2_4
Xfanout594 _04841_ vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__buf_2
X_15710_ net1350 vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__inv_2
XANTENNA__10298__A2 _04919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12922_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[16\] _03690_ net1036 vssd1
+ vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__mux2_1
X_16690_ clknet_leaf_144_wb_clk_i _02377_ _00673_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08685__C net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15641_ net1240 vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__inv_2
X_12853_ net2079 net284 net381 vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11804_ net3159 net239 net491 vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__mux2_1
X_15572_ net1400 vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__inv_2
X_12784_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] net1060 net363 _03617_
+ vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17311_ clknet_leaf_44_wb_clk_i _02998_ _01294_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14523_ net1417 vssd1 vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_25_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ _07922_ _07923_ _07925_ net613 vssd1 vssd1 vccd1 vccd1 _07926_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12708__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08663__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11612__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17242_ clknet_leaf_79_wb_clk_i _02929_ _01225_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14197__B1 net1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14454_ net1204 vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__inv_2
XANTENNA__10470__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11666_ net3145 net239 net499 vssd1 vssd1 vccd1 vccd1 _03234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12747__A1 _07588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13405_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\]
+ net596 vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__and3_1
X_10617_ net540 _06953_ _06956_ vssd1 vssd1 vccd1 vccd1 _06957_ sky130_fd_sc_hd__a21o_1
X_17173_ clknet_leaf_111_wb_clk_i _02860_ _01156_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_14385_ net1193 vssd1 vssd1 vccd1 vccd1 _00179_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11597_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] _07813_ vssd1 vssd1
+ vccd1 vccd1 _07814_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_12_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire962 _04656_ vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_12_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16124_ clknet_leaf_136_wb_clk_i _01899_ _00112_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[31\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_52_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13336_ team_01_WB.instance_to_wrap.cpu.f0.i\[14\] _07681_ net564 vssd1 vssd1 vccd1
+ vccd1 _03812_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10222__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10548_ net508 net507 net544 vssd1 vssd1 vccd1 vccd1 _06888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16055_ clknet_leaf_15_wb_clk_i _01848_ _00043_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12443__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13267_ _03756_ _03758_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[31\] net828
+ vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__14224__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10479_ _06817_ _06818_ vssd1 vssd1 vccd1 vccd1 _06819_ sky130_fd_sc_hd__and2_1
XANTENNA__09376__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15006_ net1345 vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__inv_2
X_12218_ net2888 net311 net445 vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__mux2_1
XANTENNA__09318__A _05657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13198_ net10 net837 _03738_ net3073 vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_102_Left_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12149_ net1796 net277 net452 vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__mux2_1
XANTENNA__09037__B _05338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11286__C _07111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14121__B1 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16957_ clknet_leaf_69_wb_clk_i _02644_ _00940_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11583__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15908_ net1360 vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16888_ clknet_leaf_49_wb_clk_i _02575_ _00871_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_15839_ net1330 vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09360_ _05687_ _05697_ _05698_ _05699_ vssd1 vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__or4_1
XANTENNA__13632__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08311_ net992 net965 vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_23_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17509_ clknet_leaf_50_wb_clk_i _03196_ _01492_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_111_Left_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09291_ net1009 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[22\] net910
+ vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__and3_1
XANTENNA__12618__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_126_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_13 _03663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08242_ net2928 net2714 net1048 vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1092 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_24 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_wire978_A _04635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10461__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_35 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_46 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_59_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_57 _03654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12738__A1 _07056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08173_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[108\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[100\]
+ net1044 vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_132_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10213__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10764__A3 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12353__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput120 net120 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__buf_2
Xoutput131 net131 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__buf_2
XANTENNA__08403__Y _04743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1033_A team_01_WB.instance_to_wrap.cpu.RU0.InstrRead vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xoutput142 net142 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__buf_2
XANTENNA__13163__B2 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_120_Left_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09906__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09228__A _04970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput153 net153 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
Xoutput164 net164 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__clkbuf_4
Xoutput175 net175 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__clkbuf_4
XANTENNA__11174__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout493_A _07944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16122__Q team_01_WB.instance_to_wrap.cpu.f0.data_adr\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12910__A1 _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07971__A team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14112__B1 _04259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout660_A net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout758_A _04675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_X net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09627_ _05965_ _05966_ vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout925_A net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09558_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] net626 _05897_ vssd1
+ vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__a21o_4
XTAP_TAPCELL_ROW_104_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08509_ net1079 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[18\] net925
+ vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_156_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout713_X net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10837__A net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12528__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09489_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[30\] net684 net654 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_156_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11520_ team_01_WB.instance_to_wrap.cpu.DM0.enable net717 vssd1 vssd1 vccd1 vccd1
+ _07784_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08307__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11451_ team_01_WB.instance_to_wrap.cpu.f0.i\[1\] _07671_ net325 vssd1 vssd1 vccd1
+ vccd1 _07750_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10275__C net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10402_ _06740_ _06741_ vssd1 vssd1 vccd1 vccd1 _06742_ sky130_fd_sc_hd__nand2_1
X_14170_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[6\] _04189_ net2030 vssd1
+ vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11401__A1 _07696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11382_ _07710_ vssd1 vssd1 vccd1 vccd1 _07711_ sky130_fd_sc_hd__inv_2
XANTENNA__09070__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13121_ net89 net843 net631 net1691 vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__a22o_1
X_10333_ net559 _04883_ net329 vssd1 vssd1 vccd1 vccd1 _06673_ sky130_fd_sc_hd__or3_1
XANTENNA__12263__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09358__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13052_ net2046 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[42\] net863 vssd1 vssd1
+ vccd1 vccd1 _02073_ sky130_fd_sc_hd__mux2_1
XANTENNA_input54_A wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10264_ _06221_ _06603_ _06600_ vssd1 vssd1 vccd1 vccd1 _06604_ sky130_fd_sc_hd__o21a_1
XANTENNA__14979__A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12901__A1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12003_ net2151 net242 net468 vssd1 vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__mux2_1
Xfanout1301 net1302 vssd1 vssd1 vccd1 vccd1 net1301 sky130_fd_sc_hd__buf_2
X_10195_ net1140 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[8\] net950 vssd1
+ vssd1 vccd1 vccd1 _06535_ sky130_fd_sc_hd__and3_1
X_17860_ clknet_leaf_127_wb_clk_i _03535_ _01800_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.InstrRead
+ sky130_fd_sc_hd__dfrtp_4
Xfanout1312 net1322 vssd1 vssd1 vccd1 vccd1 net1312 sky130_fd_sc_hd__clkbuf_4
Xfanout1323 net1324 vssd1 vssd1 vccd1 vccd1 net1323 sky130_fd_sc_hd__buf_4
XANTENNA__08977__A net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1334 net1344 vssd1 vssd1 vccd1 vccd1 net1334 sky130_fd_sc_hd__buf_4
XANTENNA__14103__B1 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1345 net1349 vssd1 vssd1 vccd1 vccd1 net1345 sky130_fd_sc_hd__buf_4
X_16811_ clknet_leaf_9_wb_clk_i _02498_ _00794_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1356 net1357 vssd1 vssd1 vccd1 vccd1 net1356 sky130_fd_sc_hd__buf_4
Xfanout1367 net1368 vssd1 vssd1 vccd1 vccd1 net1367 sky130_fd_sc_hd__buf_4
X_17791_ clknet_leaf_101_wb_clk_i _03467_ _01731_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[61\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_128_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout380 net382 vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__clkbuf_8
Xfanout1378 net1384 vssd1 vssd1 vccd1 vccd1 net1378 sky130_fd_sc_hd__buf_4
Xfanout1389 net1391 vssd1 vssd1 vccd1 vccd1 net1389 sky130_fd_sc_hd__buf_4
Xfanout391 net394 vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__buf_6
XANTENNA__11607__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16742_ clknet_leaf_73_wb_clk_i _02429_ _00725_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13954_ _04217_ _04219_ _04222_ vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__and3_4
XANTENNA__08122__A2_N team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12905_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[21\] _03678_ net1040 vssd1
+ vssd1 vccd1 vccd1 _03679_ sky130_fd_sc_hd__mux2_1
X_16673_ clknet_leaf_55_wb_clk_i _02360_ _00656_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13107__B net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13885_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[15\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[14\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[17\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_124_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15603__A net1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15624_ net1376 vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__inv_2
X_12836_ net2892 net218 net380 vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15555_ net1250 vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12438__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12767_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[20\] _07171_ net1032 vssd1 vssd1
+ vccd1 vccd1 _03606_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10979__A0 _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14219__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[13\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14506_ net1363 vssd1 vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__inv_2
X_11718_ _07909_ _07911_ net614 vssd1 vssd1 vccd1 vccd1 _07912_ sky130_fd_sc_hd__mux2_2
XFILLER_0_154_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15486_ net1350 vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__inv_2
X_12698_ net2941 net242 net385 vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17225_ clknet_leaf_38_wb_clk_i _02912_ _01208_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14437_ net1307 vssd1 vssd1 vccd1 vccd1 _00231_ sky130_fd_sc_hd__inv_2
XANTENNA__16207__Q net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11649_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] _07816_ vssd1 vssd1
+ vccd1 vccd1 _07857_ sky130_fd_sc_hd__xnor2_1
Xinput11 DAT_I[18] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput22 DAT_I[28] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
Xinput33 DAT_I[9] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
X_17156_ clknet_leaf_84_wb_clk_i _02843_ _01139_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput44 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_1
Xinput55 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14368_ net1208 vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__inv_2
XANTENNA__08504__X _04844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput66 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_1
Xhold806 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2341 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16107_ clknet_leaf_138_wb_clk_i _01882_ _00095_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold817 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[6\] vssd1 vssd1 vccd1 vccd1 net2352
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13319_ _07686_ _07706_ _03798_ team_01_WB.instance_to_wrap.cpu.f0.i\[18\] net587
+ vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__o221a_1
XFILLER_0_40_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold828 net138 vssd1 vssd1 vccd1 vccd1 net2363 sky130_fd_sc_hd__dlygate4sd3_1
X_17087_ clknet_leaf_41_wb_clk_i _02774_ _01070_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12173__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold839 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2374 sky130_fd_sc_hd__dlygate4sd3_1
X_14299_ net1329 vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__inv_2
XANTENNA__09349__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16038_ clknet_leaf_132_wb_clk_i net1698 _00032_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08860_ net1109 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[3\] net924 vssd1
+ vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1506 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net3041 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1517 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net3052 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_106_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_106_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08791_ net1093 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[0\] net900 vssd1
+ vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__and3_1
X_17989_ net1504 vssd1 vssd1 vccd1 vccd1 la_data_out[31] sky130_fd_sc_hd__buf_2
Xhold1528 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net3063 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_88_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1539 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net3074 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11517__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09521__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09412_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[27\] net679 net650 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[27\]
+ _05741_ vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08088__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09343_ net1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[25\] net903
+ vssd1 vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_62_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13081__A0 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12348__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout339_A _06590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09274_ _05599_ _05602_ _05612_ _05613_ vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__or4_1
XANTENNA__10434__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16117__Q team_01_WB.instance_to_wrap.cpu.f0.data_adr\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08225_ net2767 net2616 net1046 vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_151_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1150_A net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1248_A net1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09588__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08156_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[125\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[117\]
+ net1051 vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__mux2_1
XANTENNA__09884__C net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12083__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08087_ team_01_WB.instance_to_wrap.cpu.f0.i\[1\] _04524_ vssd1 vssd1 vccd1 vccd1
+ _04560_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout1036_X net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout875_A net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout496_X net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11698__A1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12811__S net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12895__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08989_ net1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[8\] net934 vssd1
+ vssd1 vccd1 vccd1 _05329_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout663_X net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09512__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout830_X net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10951_ _06468_ _06471_ vssd1 vssd1 vccd1 vccd1 _07291_ sky130_fd_sc_hd__nor2_1
XANTENNA__09124__C net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout928_X net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_123_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13670_ net1697 net568 net347 team_01_WB.instance_to_wrap.cpu.f0.i\[31\] vssd1 vssd1
+ vccd1 vccd1 _01832_ sky130_fd_sc_hd__a22o_1
X_10882_ _05566_ _06708_ vssd1 vssd1 vccd1 vccd1 _07222_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12621_ _07791_ _07945_ net574 vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08618__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15340_ net1260 vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__inv_2
X_12552_ net2144 net319 net405 vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__mux2_1
XANTENNA__10425__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11503_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[11\] _07756_ vssd1 vssd1 vccd1
+ vccd1 _07779_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15271_ net1389 vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12483_ net2072 net294 net413 vssd1 vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17010_ clknet_leaf_145_wb_clk_i _02697_ _00993_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_14222_ net3106 vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09579__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11434_ _07676_ _07685_ _07737_ _04483_ _07699_ vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__a221oi_1
XANTENNA__13375__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13089__S net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14153_ _04416_ _04436_ net604 vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11365_ team_01_WB.instance_to_wrap.cpu.f0.i\[21\] team_01_WB.instance_to_wrap.cpu.f0.i\[20\]
+ _07693_ vssd1 vssd1 vccd1 vccd1 _07694_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_4_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13104_ net63 net62 _03726_ _03727_ vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__or4_2
XFILLER_0_104_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10316_ net1129 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[18\] net948
+ vssd1 vssd1 vccd1 vccd1 _06656_ sky130_fd_sc_hd__and3_1
X_14084_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[36\] _04221_ _04259_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[20\]
+ vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__a22o_1
X_11296_ net720 net642 vssd1 vssd1 vccd1 vccd1 _07636_ sky130_fd_sc_hd__nand2_1
X_17912_ net1443 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
X_13035_ net2480 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[59\] net862 vssd1 vssd1
+ vccd1 vccd1 _02090_ sky130_fd_sc_hd__mux2_1
X_10247_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[9\] net784 net760 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[9\]
+ _06586_ vssd1 vssd1 vccd1 vccd1 _06587_ sky130_fd_sc_hd__a221o_1
Xfanout1120 net1121 vssd1 vssd1 vccd1 vccd1 net1120 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1131 net1133 vssd1 vssd1 vccd1 vccd1 net1131 sky130_fd_sc_hd__buf_2
XANTENNA__09751__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1142 net1143 vssd1 vssd1 vccd1 vccd1 net1142 sky130_fd_sc_hd__clkbuf_2
X_17843_ clknet_leaf_92_wb_clk_i net2404 _01783_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[113\]
+ sky130_fd_sc_hd__dfrtp_1
X_10178_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[10\] net740 net736 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06518_ sky130_fd_sc_hd__a22o_1
Xfanout1153 net1157 vssd1 vssd1 vccd1 vccd1 net1153 sky130_fd_sc_hd__buf_2
XANTENNA__14088__C1 net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1164 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[16\] vssd1 vssd1 vccd1 vccd1
+ net1164 sky130_fd_sc_hd__clkbuf_2
Xfanout1175 team_01_WB.instance_to_wrap.cpu.DM0.dhit vssd1 vssd1 vccd1 vccd1 net1175
+ sky130_fd_sc_hd__clkbuf_8
Xfanout1186 net1188 vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__buf_4
Xfanout1197 net1200 vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__buf_4
X_17774_ clknet_leaf_99_wb_clk_i _03450_ _01714_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[44\]
+ sky130_fd_sc_hd__dfstp_1
X_14986_ net1377 vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__inv_2
X_16725_ clknet_leaf_118_wb_clk_i _02412_ _00708_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13937_ _04227_ _04228_ vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__nand2_2
XFILLER_0_152_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13868_ net1177 net1064 net1724 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[29\]
+ sky130_fd_sc_hd__and3b_1
X_16656_ clknet_leaf_146_wb_clk_i _02343_ _00639_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12819_ net1038 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[4\] vssd1 vssd1 vccd1
+ vccd1 _03642_ sky130_fd_sc_hd__or2_2
XANTENNA__11580__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15607_ net1214 vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12168__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13799_ _04170_ _04176_ _01838_ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__a21oi_1
X_16587_ clknet_leaf_5_wb_clk_i _02274_ _00570_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13602__A2 _07553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11613__A1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15538_ net1266 vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__inv_2
XANTENNA__12810__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15469_ net1263 vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08010_ team_01_WB.instance_to_wrap.a1.WRITE_I vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__inv_2
XANTENNA__11800__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17208_ clknet_leaf_61_wb_clk_i _02895_ _01191_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold603 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2138 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmax_cap322 _07464_ vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__buf_1
XFILLER_0_142_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold614 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2149 sky130_fd_sc_hd__dlygate4sd3_1
X_17139_ clknet_leaf_17_wb_clk_i _02826_ _01122_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold625 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold636 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2171 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold647 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2182 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold658 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2193 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09990__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09961_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[3\] net785 net743 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[3\]
+ _06292_ vssd1 vssd1 vccd1 vccd1 _06301_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold669 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2204 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09209__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11129__B1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08912_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[2\] net683 _05232_ _05234_
+ _05238_ vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_55_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12631__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09892_ net1152 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[5\] net974 vssd1
+ vssd1 vccd1 vccd1 _06232_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_55_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08545__A1 net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08843_ _05163_ _05164_ _05166_ _05168_ vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__or4_1
Xhold1303 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[90\] vssd1 vssd1 vccd1 vccd1
+ net2838 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08410__A _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1314 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2849 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout191_A _07823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1325 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[112\] vssd1 vssd1 vccd1 vccd1
+ net2860 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14131__B _04396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout289_A _07941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1336 team_01_WB.instance_to_wrap.cpu.f0.num\[16\] vssd1 vssd1 vccd1 vccd1 net2871
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08774_ net598 _05110_ _05113_ vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__o21a_1
Xhold1347 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1358 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2893 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_144_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1369 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2904 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14094__A2 _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12867__A net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout456_A _07956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15243__A net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1198_A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08783__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_74_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12078__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout623_A _04628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1365_A net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09326_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[24\] net697 net685 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__a22o_1
XANTENNA__12801__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13969__Y _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09273__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11080__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09257_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[20\] net687 net667 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout411_X net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1153_X net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout509_X net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08208_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[73\] net2675 net1056 vssd1 vssd1
+ vccd1 vccd1 _03479_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09025__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09188_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[16\] net702 _05510_ _05527_
+ vssd1 vssd1 vccd1 vccd1 _05528_ sky130_fd_sc_hd__o22a_4
XANTENNA_fanout992_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08139_ _04478_ team_01_WB.instance_to_wrap.cpu.f0.num\[16\] _04497_ team_01_WB.instance_to_wrap.cpu.f0.i\[3\]
+ _04592_ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09981__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11150_ _07476_ _07489_ vssd1 vssd1 vccd1 vccd1 _07490_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout780_X net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09119__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10591__A1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout878_X net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10101_ _06438_ _06440_ vssd1 vssd1 vccd1 vccd1 _06441_ sky130_fd_sc_hd__and2_1
XANTENNA__12541__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11081_ _07420_ _07353_ vssd1 vssd1 vccd1 vccd1 _07421_ sky130_fd_sc_hd__and2b_1
XANTENNA__12868__B1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10032_ net1142 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[0\] net945 vssd1
+ vssd1 vccd1 vccd1 _06372_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_8_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09733__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11540__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14840_ net1213 vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__inv_2
XANTENNA__14085__A2 _04254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14771_ net1421 vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__inv_2
XANTENNA_input17_A DAT_I[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11983_ net1769 net303 net472 vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__mux2_1
XANTENNA__08839__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12777__A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13722_ _04108_ _04130_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[12\]
+ sky130_fd_sc_hd__nor2_1
X_16510_ clknet_leaf_5_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[8\]
+ _00493_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10934_ _05338_ net330 _07273_ net368 vssd1 vssd1 vccd1 vccd1 _07274_ sky130_fd_sc_hd__o211ai_1
X_17490_ clknet_leaf_143_wb_clk_i _03177_ _01473_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08319__X _04659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16441_ clknet_leaf_59_wb_clk_i _02195_ _00424_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13653_ _07639_ _04085_ _04086_ net728 vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__a211o_1
X_10865_ net338 _07201_ _07204_ net328 _07197_ vssd1 vssd1 vccd1 vccd1 _07205_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12604_ net2414 net261 net396 vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13596__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16372_ clknet_leaf_97_wb_clk_i _02126_ _00355_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[95\]
+ sky130_fd_sc_hd__dfrtp_1
X_13584_ _03900_ _03908_ vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__and2b_1
XANTENNA__08990__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10796_ _06036_ _07090_ vssd1 vssd1 vccd1 vccd1 _07136_ sky130_fd_sc_hd__and2_1
XANTENNA__09264__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15323_ net1253 vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12535_ net2175 net237 net403 vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10584__X _06924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12716__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15254_ net1247 vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12466_ net2475 net201 net411 vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14205_ net1556 vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__clkbuf_1
X_11417_ team_01_WB.instance_to_wrap.cpu.f0.i\[17\] _07690_ net323 vssd1 vssd1 vccd1
+ vccd1 _07732_ sky130_fd_sc_hd__o21ai_1
X_15185_ net1419 vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12397_ net2930 net206 net421 vssd1 vssd1 vccd1 vccd1 _02600_ sky130_fd_sc_hd__mux2_1
XANTENNA__08775__A1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09972__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14136_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[79\] _04235_ _04255_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[119\]
+ _04420_ vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__a221o_1
X_11348_ team_01_WB.instance_to_wrap.cpu.f0.i\[10\] team_01_WB.instance_to_wrap.cpu.f0.i\[9\]
+ net1070 vssd1 vssd1 vccd1 vccd1 _07677_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12451__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14067_ net1183 _04329_ _04355_ vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__and3_1
XANTENNA__14232__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11279_ _07042_ _07099_ _07615_ _07618_ vssd1 vssd1 vccd1 vccd1 _07619_ sky130_fd_sc_hd__a211o_1
XFILLER_0_20_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09724__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13018_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[68\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[76\]
+ net855 vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__mux2_1
XANTENNA__10334__A1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17826_ clknet_leaf_122_wb_clk_i _03502_ _01766_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[96\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14076__A2 _04241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17757_ clknet_leaf_97_wb_clk_i net2588 _01697_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_14969_ net1231 vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__inv_2
XANTENNA__11591__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10098__B1 _06436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16708_ clknet_leaf_84_wb_clk_i _02395_ _00691_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10637__A2 _06924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08490_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[23\] net680 _04795_
+ _04807_ _04816_ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__a2111o_1
X_17688_ clknet_leaf_127_wb_clk_i _03372_ _01629_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09699__C net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10919__B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15998__A net1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16639_ clknet_leaf_42_wb_clk_i _02326_ _00622_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09255__A2 _05591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09111_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[13\] net648 _05422_
+ _05430_ _05432_ vssd1 vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_45_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10935__A net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12626__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire960_A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire581_X net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09042_ net1109 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[12\] net920
+ vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14000__A2 _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold400 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1935 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold411 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1946 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout204_A _07855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold422 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1957 sky130_fd_sc_hd__dlygate4sd3_1
Xhold433 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1968 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1979 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_121_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_121_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold455 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1990 sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[15\] vssd1 vssd1 vccd1 vccd1
+ net2001 sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2012 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout902 net903 vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__buf_4
Xhold488 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2023 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09944_ _06280_ _06283_ vssd1 vssd1 vccd1 vccd1 _06284_ sky130_fd_sc_hd__and2_1
Xhold499 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2034 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout913 _04782_ vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_74_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12361__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1113_A net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout924 _04770_ vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13511__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout935 net938 vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__buf_4
XANTENNA__08778__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout946 net947 vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__clkbuf_8
X_09875_ _06209_ _06213_ _06214_ net766 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06215_ sky130_fd_sc_hd__o32a_4
XANTENNA_input9_A DAT_I[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout957 _04658_ vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__buf_6
Xhold1100 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2635 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout968 _04648_ vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__buf_4
XANTENNA_fanout194_X net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout979 net980 vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1111 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2646 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1122 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2657 sky130_fd_sc_hd__dlygate4sd3_1
X_08826_ net1104 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[1\] net884 vssd1
+ vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__and3_1
Xhold1133 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[88\] vssd1 vssd1 vccd1 vccd1
+ net2668 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1144 _02110_ vssd1 vssd1 vccd1 vccd1 net2679 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1155 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1166 team_01_WB.instance_to_wrap.cpu.f0.num\[11\] vssd1 vssd1 vccd1 vccd1 net2701
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08757_ net1099 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[4\] net898 vssd1
+ vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__and3_1
Xhold1177 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[71\] vssd1 vssd1 vccd1 vccd1
+ net2712 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout740_A net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout361_X net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1188 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[70\] vssd1 vssd1 vccd1 vccd1
+ net2723 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1199 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2734 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10089__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout838_A _03736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout459_X net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08688_ net1086 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[7\] net892 vssd1
+ vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_120_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout626_X net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10650_ net512 _06811_ net548 vssd1 vssd1 vccd1 vccd1 _06990_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09246__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09309_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[22\] net652 _05626_
+ _05640_ net705 vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__a2111o_1
X_10581_ _04710_ _06900_ vssd1 vssd1 vccd1 vccd1 _06921_ sky130_fd_sc_hd__or2_4
XANTENNA__12536__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12320_ net3052 net308 net434 vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08315__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout995_X net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10564__B _06902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12251_ net2857 net297 net442 vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11202_ _07509_ _07520_ _07531_ _07541_ vssd1 vssd1 vccd1 vccd1 _07542_ sky130_fd_sc_hd__or4_1
XANTENNA__10013__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12182_ net1945 net278 net448 vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__mux2_1
X_11133_ net541 _06924_ _07433_ _06919_ net368 vssd1 vssd1 vccd1 vccd1 _07473_ sky130_fd_sc_hd__o221a_1
XANTENNA__10580__A _04710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12271__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16990_ clknet_leaf_81_wb_clk_i _02677_ _00973_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12124__X _07957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13502__A1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08688__C net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15941_ net1418 vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__inv_2
X_11064_ _05416_ net341 vssd1 vssd1 vccd1 vccd1 _07404_ sky130_fd_sc_hd__nor2_1
XANTENNA__08914__D1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[1\] net802 net785 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06355_ sky130_fd_sc_hd__a22o_1
X_15872_ net1203 vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__inv_2
XANTENNA__14058__A2 _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17611_ clknet_leaf_129_wb_clk_i team_01_WB.instance_to_wrap.cpu.K0.next_keyvalid
+ _01552_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.keyvalid sky130_fd_sc_hd__dfrtp_4
X_14823_ net1387 vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10579__X _06919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16664__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17542_ clknet_leaf_73_wb_clk_i _03229_ _01525_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11277__C1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14754_ net1192 vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__inv_2
X_11966_ net3166 net208 net473 vssd1 vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__mux2_1
XANTENNA__09485__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13705_ team_01_WB.instance_to_wrap.cpu.c0.count\[2\] team_01_WB.instance_to_wrap.cpu.c0.count\[1\]
+ team_01_WB.instance_to_wrap.cpu.c0.count\[0\] team_01_WB.instance_to_wrap.cpu.c0.count\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__a31o_1
X_10917_ _05374_ _06591_ vssd1 vssd1 vccd1 vccd1 _07257_ sky130_fd_sc_hd__nand2_1
X_17473_ clknet_leaf_53_wb_clk_i _03160_ _01456_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_14685_ net1227 vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__inv_2
X_11897_ net3170 net213 net479 vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17919__1526 vssd1 vssd1 vccd1 vccd1 net1526 _17919__1526/LO sky130_fd_sc_hd__conb_1
XANTENNA__13569__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16424_ clknet_leaf_140_wb_clk_i _02178_ _00407_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13636_ _03862_ _03882_ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10848_ net343 _07174_ _07175_ _07187_ vssd1 vssd1 vccd1 vccd1 _07188_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_67_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09237__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12446__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13567_ _03856_ _03920_ vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__xnor2_1
X_16355_ clknet_leaf_118_wb_clk_i _02109_ _00338_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[78\]
+ sky130_fd_sc_hd__dfrtp_1
X_10779_ net530 _07118_ vssd1 vssd1 vccd1 vccd1 _07119_ sky130_fd_sc_hd__nor2_1
XANTENNA__10755__A _04844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12518_ net2523 net307 net410 vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__mux2_1
X_15306_ net1283 vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__inv_2
X_16286_ clknet_leaf_92_wb_clk_i _02040_ _00269_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13498_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[31\] net987 _03957_ _03958_
+ vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__a22o_1
X_12449_ net2416 net297 net418 vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15237_ net1286 vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13741__A1 net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15168_ net1270 vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__inv_2
XANTENNA__11752__A0 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11586__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14119_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[6\] _04249_ _04262_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[54\]
+ _04398_ vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__a221o_1
XANTENNA__12181__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15099_ net1254 vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07990_ team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1 _04488_
+ sky130_fd_sc_hd__inv_2
Xfanout209 _07847_ vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10490__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09660_ net510 _05998_ vssd1 vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__or2_1
XANTENNA__10858__A2 _06216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14049__A2 _04241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08920__A1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08611_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[11\] net906
+ net699 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[11\] vssd1 vssd1 vccd1
+ vccd1 _04951_ sky130_fd_sc_hd__a32o_1
X_17809_ clknet_leaf_121_wb_clk_i _03485_ _01749_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[79\]
+ sky130_fd_sc_hd__dfrtp_1
X_09591_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] net627 _05929_ _05930_
+ vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08542_ net1160 net620 net593 net600 vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__a211o_1
XANTENNA_clkbuf_leaf_32_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09476__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08473_ net1102 net912 vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__and2_2
XFILLER_0_58_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12356__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_832 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1063_A team_01_WB.instance_to_wrap.cpu.RU0.state\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout419_A net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09025_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[9\] net672 _05341_ _05352_
+ _05359_ vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_32_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1328_A net1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09936__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07974__A team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold230 _01978_ vssd1 vssd1 vccd1 vccd1 net1765 sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net1776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1787 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout690_A _04772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09892__C net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09400__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold263 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[11\] vssd1 vssd1 vccd1 vccd1 net1798
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_72_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold274 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1809 sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[126\] vssd1 vssd1 vccd1 vccd1
+ net1820 sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout710 net711 vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_1083 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout721 net722 vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__clkbuf_4
Xfanout732 net733 vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__clkbuf_4
X_09927_ _06257_ _06258_ _06259_ _06266_ vssd1 vssd1 vccd1 vccd1 _06267_ sky130_fd_sc_hd__or4_1
XANTENNA_clkbuf_leaf_71_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout743 net744 vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__clkbuf_8
Xfanout754 _04676_ vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout955_A _04660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout765 net766 vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__clkbuf_4
Xfanout776 _04667_ vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__clkbuf_8
Xfanout787 _04657_ vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__buf_6
X_09858_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[12\] net810 net787 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06198_ sky130_fd_sc_hd__a22o_1
Xfanout798 net799 vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__buf_6
XANTENNA__09253__X _05593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08809_ _05137_ _05140_ _05144_ _05148_ vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout743_X net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09789_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] _06128_ net623 vssd1
+ vssd1 vccd1 vccd1 _06129_ sky130_fd_sc_hd__mux2_2
X_11820_ net2250 net305 net494 vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__mux2_1
X_11751_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[1\] _07476_ net716 vssd1 vssd1
+ vccd1 vccd1 _07938_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout910_X net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09132__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08029__B net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10702_ _07039_ _07041_ net518 vssd1 vssd1 vccd1 vccd1 _07042_ sky130_fd_sc_hd__mux2_1
XANTENNA__10278__C net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14470_ net1347 vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__inv_2
X_11682_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] _07809_ vssd1 vssd1
+ vccd1 vccd1 _07883_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09219__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13421_ _03864_ _03881_ _03863_ vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__a21o_1
X_10633_ net528 _06972_ _06966_ vssd1 vssd1 vccd1 vccd1 _06973_ sky130_fd_sc_hd__o21ai_1
XANTENNA__16067__CLK clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12266__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13860__A_N net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08316__Y _04656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10234__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16140_ clknet_leaf_131_wb_clk_i _01903_ _00128_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12774__A2 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13352_ _04486_ _07678_ _03824_ vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__o21a_1
X_10564_ net555 _06902_ vssd1 vssd1 vccd1 vccd1 _06904_ sky130_fd_sc_hd__or2_2
XFILLER_0_51_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10785__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12303_ net2792 net271 net431 vssd1 vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__mux2_1
X_16071_ clknet_leaf_152_wb_clk_i _01864_ _00059_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__16035__Q team_01_WB.instance_to_wrap.cpu.f0.write_data\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13283_ _04518_ _03747_ _03770_ vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__or3_1
X_10495_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[31\] net811 vssd1 vssd1
+ vccd1 vccd1 _06835_ sky130_fd_sc_hd__and2_1
X_15022_ net1291 vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12234_ net1825 net204 net439 vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_15_Left_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08332__X _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12165_ net2254 net272 net449 vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11116_ net525 _07200_ _07455_ vssd1 vssd1 vccd1 vccd1 _07456_ sky130_fd_sc_hd__o21a_1
X_12096_ net2895 net211 net455 vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__mux2_1
X_16973_ clknet_leaf_108_wb_clk_i _02660_ _00956_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09155__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12829__A3 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11693__X _07892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11047_ net529 _06313_ vssd1 vssd1 vccd1 vccd1 _07387_ sky130_fd_sc_hd__nand2_1
X_15924_ net1360 vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__inv_2
XANTENNA__12949__B net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 DAT_I[16] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
X_15855_ net1334 vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__inv_2
X_14806_ net1261 vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_24_Left_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15786_ net1190 vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__inv_2
XANTENNA__09458__A2 _04766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12998_ net2668 net2609 net868 vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08666__A0 _04971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17525_ clknet_leaf_110_wb_clk_i _03212_ _01508_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09042__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14737_ net1196 vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__inv_2
X_11949_ net2087 net303 net476 vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_116_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_139_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17456_ clknet_leaf_109_wb_clk_i _03143_ _01439_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14668_ net1227 vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16407_ clknet_leaf_125_wb_clk_i _02161_ _00390_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12176__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13619_ _03888_ _04052_ vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17387_ clknet_leaf_10_wb_clk_i _03074_ _01370_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_14599_ net1361 vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12765__A2 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16338_ clknet_leaf_101_wb_clk_i _02092_ _00321_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[61\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_41_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16269_ clknet_leaf_156_wb_clk_i net1775 _00257_ vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_33_Left_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18008_ net635 vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09918__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09338__X _05678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13190__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07973_ team_01_WB.instance_to_wrap.cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1 _04471_
+ sky130_fd_sc_hd__inv_2
X_09712_ _06049_ _06050_ _06051_ vssd1 vssd1 vccd1 vccd1 _06052_ sky130_fd_sc_hd__or3_1
X_09643_ _05968_ _05981_ _05982_ vssd1 vssd1 vccd1 vccd1 _05983_ sky130_fd_sc_hd__or3_1
XANTENNA_clkbuf_leaf_155_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout271_A _07866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout369_A net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09574_ net1149 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[25\] net952
+ vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09449__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08525_ net1003 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[18\] net922 vssd1
+ vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__and3_1
XANTENNA__11256__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1180_A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15251__A net1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07969__A team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08456_ net1122 net1125 net1116 net1119 vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__and4b_1
XFILLER_0_148_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09887__C net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08791__C net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12086__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08387_ _04626_ _04711_ net712 vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__o21bai_1
XANTENNA_fanout703_A _04758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_154_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11003__B net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09008_ net1021 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[9\] net916 vssd1
+ vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__and3_1
XANTENNA__09909__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10280_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[19\] net730 _06617_ _06618_
+ _06619_ vssd1 vssd1 vccd1 vccd1 _06620_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_143_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout693_X net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08312__B net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17918__1525 vssd1 vssd1 vccd1 vccd1 net1525 _17918__1525/LO sky130_fd_sc_hd__conb_1
XANTENNA__09127__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout540 net541 vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout958_X net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout551 net552 vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__clkbuf_2
Xfanout562 net563 vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13872__C net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout573 _07961_ vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__clkbuf_2
X_13970_ _04218_ _04257_ vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__nor2_4
XANTENNA__09688__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout595 net596 vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__buf_2
XANTENNA__08966__C net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12921_ _05528_ net577 net360 vssd1 vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__o21ba_1
XANTENNA__12692__A1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15640_ net1209 vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__inv_2
X_12852_ net2133 net255 net382 vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11803_ net2659 net269 net491 vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__mux2_1
X_15571_ net1405 vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__inv_2
X_12783_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[15\] _07611_ net1032 vssd1 vssd1
+ vccd1 vccd1 _03617_ sky130_fd_sc_hd__mux2_1
XANTENNA__11247__A2 _07524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17310_ clknet_leaf_79_wb_clk_i _02997_ _01293_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10455__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15161__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11734_ _07798_ _07924_ vssd1 vssd1 vccd1 vccd1 _07925_ sky130_fd_sc_hd__nor2_1
X_14522_ net1366 vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_25_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08327__X _04667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09797__C net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09860__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17241_ clknet_leaf_104_wb_clk_i _02928_ _01224_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11665_ _07867_ _07869_ net611 vssd1 vssd1 vccd1 vccd1 _07870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14453_ net1224 vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__inv_2
XANTENNA__10207__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13404_ _03863_ _03864_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__nand2b_1
X_10616_ net539 _06955_ vssd1 vssd1 vccd1 vccd1 _06956_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14384_ net1193 vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__inv_2
X_17172_ clknet_leaf_66_wb_clk_i _02859_ _01155_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11596_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\]
+ _07812_ vssd1 vssd1 vccd1 vccd1 _07813_ sky130_fd_sc_hd__and3_1
XANTENNA__10758__A1 _04844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10758__B2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16123_ clknet_leaf_136_wb_clk_i _01898_ _00111_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[30\]
+ sky130_fd_sc_hd__dfrtp_4
X_13335_ _04480_ _07688_ vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__and2_1
XANTENNA__11688__X _07888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10547_ _05837_ _06829_ _06885_ net343 vssd1 vssd1 vccd1 vccd1 _06887_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_45_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08820__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap729 _04717_ vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_33_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13266_ net825 _03757_ vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__nand2_1
X_16054_ clknet_leaf_150_wb_clk_i _01847_ _00042_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\]
+ sky130_fd_sc_hd__dfrtp_4
X_10478_ _06782_ _06814_ _06815_ vssd1 vssd1 vccd1 vccd1 _06818_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11707__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12217_ net1747 net294 net446 vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__mux2_1
X_15005_ net1241 vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__inv_2
X_13197_ net11 net837 net630 net2055 vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__a22o_1
XANTENNA__08997__X _05337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11183__A1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12148_ net2784 net302 net452 vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15336__A net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16956_ clknet_leaf_50_wb_clk_i _02643_ _00939_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08997__A2_N net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12079_ net2955 net228 net459 vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__mux2_1
XANTENNA__11583__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15907_ net1367 vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_139_Right_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16887_ clknet_leaf_14_wb_clk_i _02574_ _00870_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08351__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15838_ net1330 vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__inv_2
XANTENNA__09621__X _05961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15769_ net1217 vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__inv_2
XANTENNA__11803__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08310_ net1158 net1161 net1164 net1167 vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__nor4b_1
X_17508_ clknet_leaf_82_wb_clk_i _03195_ _01491_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09290_ net1083 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[22\] net891
+ vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__and3_1
XFILLER_0_145_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10997__A1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08241_ net3068 net3026 net1049 vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__mux2_1
X_17439_ clknet_leaf_44_wb_clk_i _03126_ _01422_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_14 _04634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_25 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09500__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_36 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_47 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_58 _06098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08172_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[109\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[101\]
+ net1051 vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08811__B1 _05116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12634__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_99_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_30_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__buf_2
XFILLER_0_141_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08413__A net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput121 net121 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__buf_2
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09367__A1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput132 net132 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__buf_2
XFILLER_0_63_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13163__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput143 net143 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_28_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_140_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput154 net154 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
Xoutput165 net165 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__clkbuf_4
XANTENNA__11174__A1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1026_A net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput176 net176 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__clkbuf_4
XANTENNA__12910__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout486_A _07948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08590__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08786__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout653_A _04819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1395_A net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_67_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09626_ net511 _05964_ vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__or2_1
X_09557_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[28\] net765 _05896_ net624
+ vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__o211a_1
XANTENNA__12426__A1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout820_A _04632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout441_X net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1183_X net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout918_A _04775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08508_ net1002 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[18\] net878
+ vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09488_ _05820_ _05822_ _05827_ vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__or3_2
XFILLER_0_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09842__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_156_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08439_ net1126 net1123 net1120 net1117 vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__and4b_4
XFILLER_0_19_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout706_X net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11450_ _07673_ _07749_ vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__nor2_1
X_10401_ net371 _06739_ vssd1 vssd1 vccd1 vccd1 _06741_ sky130_fd_sc_hd__or2_1
XANTENNA__12544__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11381_ _04473_ _07709_ vssd1 vssd1 vccd1 vccd1 _07710_ sky130_fd_sc_hd__nor2_2
XFILLER_0_22_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13120_ net1675 net844 net631 team_01_WB.instance_to_wrap.a1.ADR_I\[23\] vssd1 vssd1
+ vccd1 vccd1 _02021_ sky130_fd_sc_hd__a22o_1
X_10332_ _06671_ vssd1 vssd1 vccd1 vccd1 _06672_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13154__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13051_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[35\] net2541 net862 vssd1 vssd1
+ vccd1 vccd1 _02074_ sky130_fd_sc_hd__mux2_1
X_10263_ _06533_ _06594_ _06601_ _06602_ _06499_ vssd1 vssd1 vccd1 vccd1 _06603_ sky130_fd_sc_hd__o32a_1
X_12002_ net2116 net200 net467 vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__mux2_1
XANTENNA__10291__C net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1302 net1303 vssd1 vssd1 vccd1 vccd1 net1302 sky130_fd_sc_hd__clkbuf_4
X_10194_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[8\] net804 net786 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _06534_ sky130_fd_sc_hd__a22o_1
XANTENNA_input47_A wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1313 net1315 vssd1 vssd1 vccd1 vccd1 net1313 sky130_fd_sc_hd__buf_4
Xfanout1324 net1327 vssd1 vssd1 vccd1 vccd1 net1324 sky130_fd_sc_hd__buf_4
Xfanout1335 net1337 vssd1 vssd1 vccd1 vccd1 net1335 sky130_fd_sc_hd__buf_4
X_16810_ clknet_leaf_9_wb_clk_i _02497_ _00793_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1346 net1349 vssd1 vssd1 vccd1 vccd1 net1346 sky130_fd_sc_hd__buf_4
Xfanout1357 net1362 vssd1 vssd1 vccd1 vccd1 net1357 sky130_fd_sc_hd__buf_4
X_17790_ clknet_leaf_99_wb_clk_i _03466_ _01730_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[60\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout370 _06914_ vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_128_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1368 net1369 vssd1 vssd1 vccd1 vccd1 net1368 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_128_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout381 net382 vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__clkbuf_8
Xfanout1379 net1384 vssd1 vssd1 vccd1 vccd1 net1379 sky130_fd_sc_hd__buf_4
X_16741_ clknet_leaf_51_wb_clk_i _02428_ _00724_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout392 net394 vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__buf_8
XFILLER_0_89_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13953_ _04217_ _04220_ _04228_ vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__and3_4
X_12904_ _05591_ net577 net360 vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__o21ba_1
X_16672_ clknet_leaf_48_wb_clk_i _02359_ _00655_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13884_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[13\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[12\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[11\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__or4bb_1
XANTENNA__13107__C net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10140__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15623_ net1389 vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12835_ net3054 net221 net379 vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12719__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11623__S net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10428__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15554_ net1319 vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12766_ net1815 net639 net607 _03605_ vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09833__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10979__A1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14505_ net1364 vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__inv_2
X_11717_ _07801_ _07910_ vssd1 vssd1 vccd1 vccd1 _07911_ sky130_fd_sc_hd__nor2_1
X_15485_ net1236 vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__inv_2
X_12697_ net2670 net201 net383 vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17224_ clknet_leaf_64_wb_clk_i _02911_ _01207_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11648_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[22\] _07154_ net713 vssd1 vssd1
+ vccd1 vccd1 _07856_ sky130_fd_sc_hd__mux2_1
X_14436_ net1228 vssd1 vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput12 DAT_I[19] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
Xinput23 DAT_I[29] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput34 gpio_in[16] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_1
Xinput45 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_1
X_17155_ clknet_leaf_22_wb_clk_i _02842_ _01138_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11579_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[31\] _06961_ net715 vssd1 vssd1
+ vccd1 vccd1 _07796_ sky130_fd_sc_hd__mux2_1
X_14367_ net1208 vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__inv_2
XANTENNA__12454__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput56 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput67 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11211__X _07551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold807 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2342 sky130_fd_sc_hd__dlygate4sd3_1
X_16106_ clknet_leaf_138_wb_clk_i _01881_ _00094_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[13\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold818 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2353 sky130_fd_sc_hd__dlygate4sd3_1
X_13318_ team_01_WB.instance_to_wrap.cpu.f0.i\[17\] net610 _07703_ vssd1 vssd1 vccd1
+ vccd1 _03798_ sky130_fd_sc_hd__and3_1
X_17086_ clknet_leaf_82_wb_clk_i _02773_ _01069_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold829 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2364 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14298_ net1329 vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__inv_2
XANTENNA__13145__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16037_ clknet_leaf_133_wb_clk_i _01831_ _00031_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13249_ net2716 net355 net351 team_01_WB.instance_to_wrap.cpu.f0.i\[1\] vssd1 vssd1
+ vccd1 vccd1 _01901_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11594__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08572__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08790_ net1094 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[0\] net929 vssd1
+ vssd1 vccd1 vccd1 _05130_ sky130_fd_sc_hd__and3_1
XANTENNA__10702__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1507 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net3042 sky130_fd_sc_hd__dlygate4sd3_1
X_17988_ net1503 vssd1 vssd1 vccd1 vccd1 la_data_out[30] sky130_fd_sc_hd__buf_2
Xhold1518 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net3053 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1529 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net3064 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_88_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09064__A net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16939_ clknet_leaf_9_wb_clk_i _02626_ _00922_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_146_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_146_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09411_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[27\] net683 _05750_
+ net705 vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__a211o_1
XFILLER_0_95_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12629__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09342_ _05681_ vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08408__A _04738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09273_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[20\] net650 net648 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[20\]
+ _05598_ vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17917__1524 vssd1 vssd1 vccd1 vccd1 net1524 _17917__1524/LO sky130_fd_sc_hd__conb_1
XFILLER_0_145_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout234_A net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10376__C net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08224_ net2529 net2381 net1056 vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14030__B1 _04236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08155_ net1820 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[118\] net1044 vssd1 vssd1
+ vccd1 vccd1 _03532_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout401_A _03566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12364__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10817__S1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1143_A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08414__Y _04754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08086_ _04529_ _04539_ _04558_ vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__o21bai_1
XANTENNA__13136__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10960__X _07300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1310_A net1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11147__A1 _06906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1408_A net1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout770_A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12895__A1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout391_X net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08430__X _04770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout489_X net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14097__B1 _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08988_ net1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[8\] net939 vssd1
+ vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_106_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout656_X net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10658__A0 _06216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11791__X _07944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1398_X net1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10950_ net562 _07189_ _07270_ _07289_ vssd1 vssd1 vccd1 vccd1 _07290_ sky130_fd_sc_hd__a31o_2
XANTENNA__15704__A net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10122__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09609_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[24\] net783 net773 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__a22o_1
XANTENNA__09702__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout823_X net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10881_ _05566_ net330 _07220_ vssd1 vssd1 vccd1 vccd1 _07221_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12539__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12620_ net2017 net291 net396 vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__mux2_1
XANTENNA__09815__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12551_ net1984 net305 net405 vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11502_ net1666 net876 _07758_ _07778_ vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__o22a_1
X_12482_ net2466 net296 net414 vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__mux2_1
X_15270_ net1381 vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__inv_2
XANTENNA__14021__B1 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11433_ _07678_ _07701_ _07741_ net324 vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__o211a_1
X_14221_ net1593 vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12274__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14055__A _04230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14152_ _04222_ _04228_ _04237_ _04289_ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__a31o_1
X_11364_ team_01_WB.instance_to_wrap.cpu.f0.i\[19\] _07692_ vssd1 vssd1 vccd1 vccd1
+ _07693_ sky130_fd_sc_hd__and2_1
X_13103_ net59 net60 vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__nand2_1
XANTENNA__13127__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10315_ net990 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[18\] net975 vssd1
+ vssd1 vccd1 vccd1 _06655_ sky130_fd_sc_hd__and3_1
X_14083_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[60\] _04260_ _04261_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[116\]
+ _04370_ vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__a221o_1
X_11295_ net725 _04838_ vssd1 vssd1 vccd1 vccd1 _07635_ sky130_fd_sc_hd__nor2_1
X_17911_ net1442 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
X_13034_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[52\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[60\]
+ net855 vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__mux2_1
X_10246_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[9\] net790 _06584_ _06585_
+ vssd1 vssd1 vccd1 vccd1 _06586_ sky130_fd_sc_hd__a211o_1
XANTENNA__08340__X _04680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12886__A1 _05726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1110 net1113 vssd1 vssd1 vccd1 vccd1 net1110 sky130_fd_sc_hd__clkbuf_2
Xfanout1121 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[22\] vssd1 vssd1 vccd1 vccd1
+ net1121 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11618__S net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1132 net1133 vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__clkbuf_2
X_17842_ clknet_leaf_122_wb_clk_i net2861 _01782_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[112\]
+ sky130_fd_sc_hd__dfrtp_1
X_10177_ _06505_ _06508_ _06513_ _06516_ vssd1 vssd1 vccd1 vccd1 _06517_ sky130_fd_sc_hd__nor4_1
Xfanout1143 net1144 vssd1 vssd1 vccd1 vccd1 net1143 sky130_fd_sc_hd__buf_2
Xfanout1154 net1156 vssd1 vssd1 vccd1 vccd1 net1154 sky130_fd_sc_hd__clkbuf_2
Xfanout1165 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[16\] vssd1 vssd1 vccd1 vccd1
+ net1165 sky130_fd_sc_hd__clkbuf_2
Xfanout1176 team_01_WB.instance_to_wrap.cpu.f0.state\[4\] vssd1 vssd1 vccd1 vccd1
+ net1176 sky130_fd_sc_hd__buf_2
X_17773_ clknet_leaf_95_wb_clk_i _03449_ _01713_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[43\]
+ sky130_fd_sc_hd__dfrtp_1
X_14985_ net1294 vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__inv_2
Xfanout1187 net1188 vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__clkbuf_2
Xfanout1198 net1200 vssd1 vssd1 vccd1 vccd1 net1198 sky130_fd_sc_hd__buf_4
XFILLER_0_135_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10649__A0 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16724_ clknet_leaf_22_wb_clk_i _02411_ _00707_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13936_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[3\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__nor2_2
XFILLER_0_53_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16655_ clknet_leaf_35_wb_clk_i _02342_ _00638_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12449__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13867_ net1177 net1064 net1668 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[28\]
+ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_83_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15606_ net1256 vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__inv_2
X_12818_ net1035 _07449_ vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__nand2_1
XANTENNA__11580__C team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16586_ clknet_leaf_5_wb_clk_i _02273_ _00569_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09267__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13798_ _04159_ _04174_ _04179_ _04154_ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__a22o_1
XANTENNA__09806__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15537_ net1393 vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09050__C net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11613__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12749_ net1838 net640 net608 _03593_ vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12810__B2 _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10196__C net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15468_ net1257 vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__inv_2
XANTENNA__14012__B1 _04244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17207_ clknet_leaf_13_wb_clk_i _02894_ _01190_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_14419_ net1308 vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_7_Left_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12184__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15399_ net1395 vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold604 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2139 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13771__C1 net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17138_ clknet_leaf_144_wb_clk_i _02825_ _01121_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold615 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 net2150
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2161 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold637 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2172 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13118__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold648 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2183 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold659 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2194 sky130_fd_sc_hd__dlygate4sd3_1
X_09960_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[3\] net747 net735 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06300_ sky130_fd_sc_hd__a22o_1
X_17069_ clknet_leaf_108_wb_clk_i _02756_ _01052_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13523__C1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08911_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[2\] net681 _05230_ _05236_
+ _05240_ vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__a2111o_1
X_09891_ net1153 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[5\] net950 vssd1
+ vssd1 vccd1 vccd1 _06231_ sky130_fd_sc_hd__and3_1
XANTENNA__12877__A1 _05802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08842_ _05179_ _05180_ _05181_ vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__or3_1
Xhold1304 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[17\] vssd1 vssd1 vccd1 vccd1
+ net2839 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14079__B1 _04245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10352__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08410__B net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1315 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[111\] vssd1 vssd1 vccd1 vccd1
+ net2850 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1326 _03518_ vssd1 vssd1 vccd1 vccd1 net2861 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08773_ net603 _05112_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__or2_1
Xhold1337 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[102\] vssd1 vssd1 vccd1 vccd1
+ net2872 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1348 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[15\] vssd1 vssd1 vccd1 vccd1
+ net2883 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1359 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[63\] vssd1 vssd1 vccd1 vccd1
+ net2894 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_144_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12867__B _07756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12359__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1093_A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout449_A _07958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09258__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09325_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[24\] net678 net671 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[24\]
+ _05663_ vssd1 vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__a221o_1
XANTENNA__12801__A1 _07269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1260_A net1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09256_ net1080 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[20\] net935
+ vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14003__B1 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08207_ net2359 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[66\] net1052 vssd1 vssd1
+ vccd1 vccd1 _03480_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_43_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_133_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09187_ _05514_ _05518_ _05522_ _05526_ vssd1 vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__or4_1
XANTENNA__12094__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout404_X net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08138_ _04478_ team_01_WB.instance_to_wrap.cpu.f0.num\[16\] team_01_WB.instance_to_wrap.cpu.f0.num\[10\]
+ _04483_ _04591_ vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__o221ai_1
XTAP_TAPCELL_ROW_79_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09430__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout985_A _04629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08784__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11011__B net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08304__C net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08069_ _04542_ _04543_ _04544_ _04545_ vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__or4_1
X_10100_ _05043_ _06439_ vssd1 vssd1 vccd1 vccd1 _06440_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11080_ _05618_ net507 _07355_ net508 _05594_ vssd1 vssd1 vccd1 vccd1 _07420_ sky130_fd_sc_hd__o32a_1
XANTENNA_fanout773_X net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10031_ net1142 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[0\] net951 vssd1
+ vssd1 vccd1 vccd1 _06371_ sky130_fd_sc_hd__and3_1
XANTENNA__08536__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11540__B2 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout940_X net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09135__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14770_ net1286 vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11982_ net2187 net280 net472 vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__mux2_1
XANTENNA__12777__B team_01_WB.instance_to_wrap.cpu.f0.data_adr\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08974__C net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13721_ net2896 _04107_ vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__nor2_1
X_10933_ _06919_ _06912_ _07272_ vssd1 vssd1 vccd1 vccd1 _07273_ sky130_fd_sc_hd__mux2_1
XANTENNA__12269__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16440_ clknet_leaf_75_wb_clk_i _02194_ _00423_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10864_ _07118_ _07200_ net525 vssd1 vssd1 vccd1 vccd1 _07204_ sky130_fd_sc_hd__mux2_1
X_13652_ net198 net194 _07930_ net645 vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__o211a_1
XANTENNA__09249__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13889__A net1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12603_ net2208 net267 net395 vssd1 vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16371_ clknet_leaf_119_wb_clk_i _02125_ _00354_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[94\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13583_ net988 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] _04027_ _04028_
+ vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__a22o_1
X_10795_ net562 _07115_ _07116_ _07134_ vssd1 vssd1 vccd1 vccd1 _07135_ sky130_fd_sc_hd__a31o_2
XFILLER_0_26_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11901__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15322_ net1371 vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12534_ net2795 net269 net403 vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08335__X _04675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15253_ net1276 vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__inv_2
X_12465_ net3135 net204 net411 vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__mux2_1
X_14204_ net2507 vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11416_ _07692_ net323 _07730_ vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__and3b_1
X_12396_ net3027 net247 net421 vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__mux2_1
XANTENNA__09421__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15184_ net1276 vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11347_ team_01_WB.instance_to_wrap.cpu.f0.i\[6\] _07675_ vssd1 vssd1 vccd1 vccd1
+ _07676_ sky130_fd_sc_hd__and2_1
XANTENNA__08775__A2 _05110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09972__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14135_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[87\] _04251_ _04268_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[79\]
+ vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_728 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09607__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11278_ _05595_ net508 _07616_ _07617_ vssd1 vssd1 vccd1 vccd1 _07618_ sky130_fd_sc_hd__o22a_1
X_14066_ _04332_ _04341_ _04348_ _04354_ vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__or4_1
X_10229_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[9\] net776 net752 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06569_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_33_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13017_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[69\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[77\]
+ net864 vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17916__1523 vssd1 vssd1 vccd1 vccd1 net1523 _17916__1523/LO sky130_fd_sc_hd__conb_1
XANTENNA__11531__B2 net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17825_ clknet_leaf_121_wb_clk_i net2641 _01765_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[95\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1 team_01_WB.instance_to_wrap.cpu.K0.state vssd1 vssd1 vccd1 vccd1 net1536 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09045__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17756_ clknet_leaf_92_wb_clk_i _03432_ _01696_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_22_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14968_ net1213 vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__inv_2
XANTENNA__10098__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11591__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16707_ clknet_leaf_29_wb_clk_i _02394_ _00690_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13919_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[12\] _04212_ _04213_ vssd1
+ vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__o21a_1
XANTENNA__12179__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17687_ clknet_leaf_127_wb_clk_i _03371_ _01628_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_14899_ net1392 vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__inv_2
X_16638_ clknet_leaf_81_wb_clk_i _02325_ _00621_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16569_ clknet_leaf_104_wb_clk_i _02256_ _00552_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09110_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[13\] net683 _05421_
+ _05442_ net708 vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11811__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12795__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09041_ net1169 net620 net593 vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__a21o_1
XFILLER_0_26_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold401 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net1936 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09412__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_83 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold412 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1947 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold423 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1958 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold434 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1969 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08766__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold445 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1980 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12642__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1026 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold456 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net1991 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold467 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2002 sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2013 sky130_fd_sc_hd__dlygate4sd3_1
Xhold489 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2024 sky130_fd_sc_hd__dlygate4sd3_1
X_09943_ net554 _06282_ vssd1 vssd1 vccd1 vccd1 _06283_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_74_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_61_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout903 _04788_ vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__buf_4
XANTENNA__08421__A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10670__B _06398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout914 _04779_ vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__buf_4
XFILLER_0_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10493__A_N net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout925 net928 vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_146_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout936 net938 vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__buf_4
XANTENNA_fanout399_A _03566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_wb_clk_i_X clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13511__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09874_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[12\] net750 net747 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[12\]
+ _06197_ vssd1 vssd1 vccd1 vccd1 _06214_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_5_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout958 net962 vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__buf_4
XANTENNA__11522__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1101 team_01_WB.instance_to_wrap.cpu.f0.num\[13\] vssd1 vssd1 vccd1 vccd1 net2636
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout969 _04648_ vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1106_A net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1112 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[24\] vssd1 vssd1 vccd1 vccd1
+ net2647 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1123 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2658 sky130_fd_sc_hd__dlygate4sd3_1
X_08825_ net1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[1\] net913 vssd1
+ vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__and3_1
Xhold1134 team_01_WB.instance_to_wrap.cpu.f0.num\[30\] vssd1 vssd1 vccd1 vccd1 net2669
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1145 team_01_WB.instance_to_wrap.cpu.f0.num\[19\] vssd1 vssd1 vccd1 vccd1 net2680
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout187_X net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1156 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2691 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15254__A net1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1167 team_01_WB.instance_to_wrap.cpu.f0.num\[4\] vssd1 vssd1 vccd1 vccd1 net2702
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08756_ net1017 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[4\] net927 vssd1
+ vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__and3_1
XANTENNA__13275__A1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1178 _03477_ vssd1 vssd1 vccd1 vccd1 net2713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1189 _03476_ vssd1 vssd1 vccd1 vccd1 net2724 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08794__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12089__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08687_ net1085 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[7\] net944 vssd1
+ vssd1 vccd1 vccd1 _05027_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_120_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1096_X net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout900_A net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10941__A1_N net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09308_ _05644_ _05645_ _05646_ _05647_ vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10580_ _04710_ _06900_ vssd1 vssd1 vccd1 vccd1 _06920_ sky130_fd_sc_hd__nor2_4
XANTENNA__09651__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10261__A1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09239_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[21\] net687 net666 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1430_X net1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12250_ net2575 net276 net440 vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout890_X net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09403__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout988_X net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11201_ _07533_ _07539_ _07540_ vssd1 vssd1 vccd1 vccd1 _07541_ sky130_fd_sc_hd__or3_2
XFILLER_0_31_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12181_ net2110 net301 net448 vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12552__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11761__A1 _07831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11132_ net337 _07433_ vssd1 vssd1 vccd1 vccd1 _07472_ sky130_fd_sc_hd__nand2_1
XANTENNA__08969__C net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold990 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2525 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_79_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13502__A2 _07019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11063_ _07379_ _07402_ vssd1 vssd1 vccd1 vccd1 _07403_ sky130_fd_sc_hd__nand2_1
X_15940_ net1361 vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__inv_2
XANTENNA__11513__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10014_ _06350_ _06351_ _06352_ _06353_ vssd1 vssd1 vccd1 vccd1 _06354_ sky130_fd_sc_hd__or4_1
XANTENNA__09182__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15871_ net1203 vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__inv_2
X_17610_ clknet_leaf_129_wb_clk_i team_01_WB.instance_to_wrap.cpu.K0.next_state _01551_
+ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.state sky130_fd_sc_hd__dfrtp_1
X_14822_ net1404 vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__inv_2
X_17541_ clknet_leaf_47_wb_clk_i _03228_ _01524_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_14753_ net1188 vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11965_ net2852 net245 net473 vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13704_ net2868 _04101_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[4\]
+ sky130_fd_sc_hd__xor2_1
X_17472_ clknet_leaf_46_wb_clk_i _03159_ _01455_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10916_ _07254_ _07255_ net521 vssd1 vssd1 vccd1 vccd1 _07256_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14684_ net1306 vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__inv_2
XANTENNA__10101__A _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_106_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11896_ net2370 net214 net479 vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_88_Left_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16423_ clknet_leaf_141_wb_clk_i _02177_ _00406_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13635_ net987 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] _04071_ _04072_
+ vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__a22o_1
X_10847_ net558 _07186_ _07184_ vssd1 vssd1 vccd1 vccd1 _07187_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_73_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11631__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16354_ clknet_leaf_101_wb_clk_i _02108_ _00337_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[77\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_137_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13566_ net986 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] _04013_ _04014_
+ vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__a22o_1
X_10778_ _07104_ _07117_ net514 vssd1 vssd1 vccd1 vccd1 _07118_ sky130_fd_sc_hd__mux2_1
XANTENNA__08506__A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10755__B net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15305_ net1293 vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__inv_2
XANTENNA__10252__A1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12517_ net1921 net310 net408 vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16285_ clknet_leaf_123_wb_clk_i _02039_ _00268_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13497_ net721 _06961_ net1074 vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15236_ net1220 vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__inv_2
X_12448_ net1980 net278 net416 vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15167_ net1318 vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__inv_2
XANTENNA__12462__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12379_ net1959 net252 net425 vssd1 vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_97_Left_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14118_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[46\] _04246_ _04250_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[126\]
+ _04403_ vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__a221o_1
XANTENNA__11586__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15098_ net1370 vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14151__C1 net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14049_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[91\] _04241_ _04258_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[59\]
+ _04337_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10858__A3 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_145_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_4__f_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11806__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08920__A2 _05258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08610_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[11\] net687 net652 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__a22o_1
X_09590_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[25\] net765 net624 vssd1
+ vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__o21a_1
X_17808_ clknet_leaf_120_wb_clk_i _03484_ _01748_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[78\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17739_ clknet_leaf_92_wb_clk_i _03415_ _01679_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_08541_ net592 net591 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[18\] net701
+ vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__o2bb2a_4
XANTENNA__09503__C net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08472_ net1081 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[23\] net878
+ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__and3_1
XANTENNA__09527__A1_N net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_947 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12637__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12768__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_139_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10665__B _06280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08987__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13980__A2 _04236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09024_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[9\] net669 _05345_ _05351_
+ _05354_ vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout1056_A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13193__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold220 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1755 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12372__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold231 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1766 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12225__X _07962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold242 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1777 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1223_A net1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold253 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[123\] vssd1 vssd1 vccd1 vccd1
+ net1788 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1799 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08789__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold275 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[10\] vssd1 vssd1 vccd1 vccd1
+ net1810 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout700 _04760_ vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__buf_4
Xhold286 _03532_ vssd1 vssd1 vccd1 vccd1 net1821 sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1832 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout711 _04728_ vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__clkbuf_4
X_09926_ _06260_ _06261_ _06265_ vssd1 vssd1 vccd1 vccd1 _06266_ sky130_fd_sc_hd__or3_1
XFILLER_0_102_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout722 _04721_ vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__buf_2
XFILLER_0_141_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout733 _04688_ vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__buf_4
XANTENNA__13496__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout744 _04684_ vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__buf_4
Xfanout755 _04675_ vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07990__A team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout766 net767 vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__buf_4
Xfanout777 _04666_ vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__clkbuf_8
X_09857_ net1156 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[12\] net971
+ vssd1 vssd1 vccd1 vccd1 _06197_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout850_A net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout788 _04657_ vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout471_X net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout799 _04649_ vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__buf_6
XANTENNA_fanout569_X net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout948_A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08911__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08808_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[0\] net684 _05145_ _05146_
+ _05147_ vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13248__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09788_ _06111_ _06118_ _06126_ _06127_ vssd1 vssd1 vccd1 vccd1 _06128_ sky130_fd_sc_hd__o31a_2
X_08739_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[4\] net936 vssd1
+ vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout736_X net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15712__A net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11750_ net2341 net317 net501 vssd1 vssd1 vccd1 vccd1 _03217_ sky130_fd_sc_hd__mux2_1
XANTENNA__09872__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10701_ _07040_ vssd1 vssd1 vccd1 vccd1 _07041_ sky130_fd_sc_hd__inv_2
XANTENNA__12547__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11681_ net719 _07611_ net615 _07881_ vssd1 vssd1 vccd1 vccd1 _07882_ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout903_X net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12759__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13420_ _03867_ _03880_ _03866_ vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__a21o_1
X_10632_ net514 _06969_ _06970_ _06971_ vssd1 vssd1 vccd1 vccd1 _06972_ sky130_fd_sc_hd__a31o_1
XFILLER_0_153_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08326__A net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17915__1522 vssd1 vssd1 vccd1 vccd1 net1522 _17915__1522/LO sky130_fd_sc_hd__conb_1
X_10563_ net555 _06902_ vssd1 vssd1 vccd1 vccd1 _06903_ sky130_fd_sc_hd__nor2_2
X_13351_ team_01_WB.instance_to_wrap.cpu.f0.i\[11\] net610 vssd1 vssd1 vccd1 vccd1
+ _03824_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10785__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12302_ net2932 net243 net433 vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__mux2_1
X_16070_ clknet_leaf_154_wb_clk_i _01863_ _00058_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\]
+ sky130_fd_sc_hd__dfstp_4
XFILLER_0_133_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13282_ team_01_WB.instance_to_wrap.cpu.f0.i\[24\] _03746_ team_01_WB.instance_to_wrap.cpu.f0.i\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__a21oi_1
X_10494_ net1130 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[31\] net984
+ vssd1 vssd1 vccd1 vccd1 _06834_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15021_ net1266 vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__inv_2
XANTENNA__13184__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11687__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12282__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12233_ net2827 net272 net441 vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__mux2_1
XANTENNA__10537__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09157__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12164_ net2619 net209 net449 vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11115_ _06905_ _07303_ _07454_ _05263_ vssd1 vssd1 vccd1 vccd1 _07455_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__16051__Q team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16972_ clknet_leaf_19_wb_clk_i _02659_ _00955_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_12095_ net2920 net214 net457 vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__mux2_1
X_11046_ net529 _06313_ vssd1 vssd1 vccd1 vccd1 _07386_ sky130_fd_sc_hd__or2_1
X_15923_ net1367 vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11626__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15854_ net1334 vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__inv_2
XANTENNA__10170__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13239__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14805_ net1287 vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__inv_2
X_15785_ net1190 vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__inv_2
X_12997_ net2935 net2745 net866 vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17524_ clknet_leaf_66_wb_clk_i _03211_ _01507_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_14736_ net1196 vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11948_ net1884 net280 net476 vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__mux2_1
XANTENNA__08666__A1 _05005_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09863__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17455_ clknet_leaf_37_wb_clk_i _03142_ _01438_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_14667_ net1228 vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__inv_2
XANTENNA__12457__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11879_ net2508 net285 net485 vssd1 vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__mux2_1
X_16406_ clknet_leaf_124_wb_clk_i _02160_ _00389_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13618_ net987 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] _04057_ _04058_
+ vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17386_ clknet_leaf_30_wb_clk_i _03073_ _01369_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_14598_ net1360 vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16337_ clknet_leaf_118_wb_clk_i _02091_ _00320_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[60\]
+ sky130_fd_sc_hd__dfstp_1
X_13549_ net986 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] _03999_ _04000_
+ vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11973__A1 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16268_ clknet_leaf_153_wb_clk_i net1716 _00256_ vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__dfrtp_1
X_18007_ net637 vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15219_ net1421 vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11597__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12192__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16199_ clknet_leaf_159_wb_clk_i _01959_ _00187_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10528__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07972_ team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1 _04470_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_96_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09711_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[21\] net761 net743 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__a22o_1
XANTENNA__08354__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09642_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[23\] net807 _05972_
+ _05974_ _05980_ vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_78_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09573_ net1149 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[25\] net946
+ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__and3_1
XANTENNA__08106__B1 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout264_A _07880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08524_ net1001 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[18\] net901
+ vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__and3_1
XANTENNA__13650__A1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09530__A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12367__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08455_ net1001 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[23\] net897 vssd1
+ vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout431_A _07964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout529_A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08386_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[6\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[2\]
+ _04623_ _04725_ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__nor4_1
XFILLER_0_92_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1059_X net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08433__X _04773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout898_A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13166__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09007_ net1100 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[9\] net884 vssd1
+ vssd1 vccd1 vccd1 _05347_ sky130_fd_sc_hd__and3_1
XFILLER_0_143_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09909__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[5\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11177__C1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1226_X net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10519__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09385__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout686_X net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout530 net532 vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__clkbuf_4
Xfanout541 net542 vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__clkbuf_4
Xfanout552 _05151_ vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__buf_2
X_09909_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[5\] net765 net624 vssd1
+ vssd1 vccd1 vccd1 _06249_ sky130_fd_sc_hd__o21a_1
XANTENNA__14130__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09705__A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout563 _04747_ vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout853_X net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout574 _07961_ vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__buf_1
X_12920_ net359 _03688_ _03689_ net872 net1563 vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__a32o_1
Xfanout596 _04840_ vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10152__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12851_ net1978 net257 net381 vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_9__f_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_9__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__10289__C net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11802_ net2452 net242 net493 vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15570_ net1290 vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_4_3__f_wb_clk_i_X clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12782_ net2053 net640 net608 _03616_ vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08982__C net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14521_ net1364 vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11733_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] _07797_ vssd1 vssd1 vccd1
+ vccd1 _07924_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12277__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17240_ clknet_leaf_38_wb_clk_i _02927_ _01223_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14452_ net1204 vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__inv_2
X_11664_ _07813_ _07868_ vssd1 vssd1 vccd1 vccd1 _07869_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13403_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] net595 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10615_ net547 _06366_ _06399_ vssd1 vssd1 vccd1 vccd1 _06955_ sky130_fd_sc_hd__o21ai_1
X_17171_ clknet_leaf_17_wb_clk_i _02858_ _01154_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_148_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14383_ net1195 vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11595_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\]
+ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] _07809_ vssd1 vssd1 vccd1 vccd1
+ _07812_ sky130_fd_sc_hd__and4_1
XANTENNA__10758__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16122_ clknet_leaf_136_wb_clk_i _01897_ _00110_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13334_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[17\] net828 _03809_ _03810_
+ vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_12_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09439__X _05779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10546_ _05837_ _06829_ _06885_ vssd1 vssd1 vccd1 vccd1 _06886_ sky130_fd_sc_hd__a21o_1
XANTENNA__13157__B1 _03734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16053_ clknet_leaf_4_wb_clk_i _01846_ _00041_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_13265_ _04518_ _03750_ _03755_ _04621_ _04466_ vssd1 vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_110_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10477_ net512 _05933_ _06816_ vssd1 vssd1 vccd1 vccd1 _06817_ sky130_fd_sc_hd__o21ai_2
XANTENNA__11707__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15004_ net1246 vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12216_ net2230 net296 net446 vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__mux2_1
XANTENNA__09376__A2 _04776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13196_ net12 net837 net630 net2132 vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12147_ net2177 net282 net454 vssd1 vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__mux2_1
XANTENNA__10391__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14121__A2 _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12078_ net2782 net285 net462 vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__mux2_1
X_16955_ clknet_leaf_70_wb_clk_i _02642_ _00938_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11029_ _05455_ net373 vssd1 vssd1 vccd1 vccd1 _07369_ sky130_fd_sc_hd__nor2_1
X_15906_ net1352 vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16886_ clknet_leaf_12_wb_clk_i _02573_ _00869_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10143__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15837_ net1331 vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__inv_2
XANTENNA__09053__C net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10199__C net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15768_ net1199 vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__inv_2
XANTENNA__09836__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08892__C net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14719_ net1189 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__inv_2
X_17507_ clknet_leaf_25_wb_clk_i _03194_ _01490_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12187__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15699_ net1419 vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__inv_2
XANTENNA__10496__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08240_ net2400 net2321 net1057 vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17438_ clknet_leaf_85_wb_clk_i _03125_ _01421_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_15 _07289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_37 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_48 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08171_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[110\] net2872 net1043 vssd1 vssd1
+ vccd1 vccd1 _03516_ sky130_fd_sc_hd__mux2_1
X_17369_ clknet_leaf_102_wb_clk_i _03056_ _01352_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_59 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08811__A1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13148__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__buf_2
XFILLER_0_24_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__buf_2
Xoutput122 net122 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__buf_2
XFILLER_0_141_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09367__A2 _05705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput133 net133 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__buf_2
XFILLER_0_101_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput144 net144 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__buf_2
XFILLER_0_2_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput155 net155 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
XFILLER_0_100_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput166 net166 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__clkbuf_4
XANTENNA__12371__A1 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput177 net177 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_56_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12650__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08700__Y _05040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10382__B1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1019_A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14112__A2 _04230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_68_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout381_A net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout479_A _07949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09625_ net511 _05964_ vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_67_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout646_A _04825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09556_ _05888_ _05889_ _05893_ _05895_ vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__or4_1
XANTENNA__09827__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13623__A1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08507_ net1160 net620 net593 vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__a21o_1
XANTENNA__11634__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12097__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout813_A net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout434_X net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09487_ _05823_ _05824_ _05825_ _05826_ vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_156_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08438_ net1016 net938 vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_156_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08307__C net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11014__B net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08369_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] net1169 vssd1 vssd1 vccd1
+ vccd1 _04709_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout601_X net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10400_ net371 _06739_ vssd1 vssd1 vccd1 vccd1 _06740_ sky130_fd_sc_hd__nand2_2
XFILLER_0_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11380_ team_01_WB.instance_to_wrap.cpu.f0.i\[20\] _07707_ vssd1 vssd1 vccd1 vccd1
+ _07709_ sky130_fd_sc_hd__nand2_2
XANTENNA__13139__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10331_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] net625 _06669_ _06670_
+ vssd1 vssd1 vccd1 vccd1 _06671_ sky130_fd_sc_hd__a22o_4
XANTENNA__08323__B net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10262_ _06500_ _06530_ vssd1 vssd1 vccd1 vccd1 _06602_ sky130_fd_sc_hd__nor2_1
XANTENNA__09358__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13050_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[36\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[44\]
+ net858 vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout970_X net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09138__C net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12001_ net1830 net204 net467 vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__mux2_1
X_10193_ _06499_ _06500_ _06532_ vssd1 vssd1 vccd1 vccd1 _06533_ sky130_fd_sc_hd__or3_1
XANTENNA__12560__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1303 net1304 vssd1 vssd1 vccd1 vccd1 net1303 sky130_fd_sc_hd__clkbuf_4
Xfanout1314 net1315 vssd1 vssd1 vccd1 vccd1 net1314 sky130_fd_sc_hd__buf_4
Xfanout1325 net1327 vssd1 vssd1 vccd1 vccd1 net1325 sky130_fd_sc_hd__buf_4
XANTENNA__08977__C net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14103__A2 _04246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1336 net1337 vssd1 vssd1 vccd1 vccd1 net1336 sky130_fd_sc_hd__buf_4
Xfanout1347 net1348 vssd1 vssd1 vccd1 vccd1 net1347 sky130_fd_sc_hd__buf_4
Xfanout360 net361 vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__buf_2
Xfanout1358 net1362 vssd1 vssd1 vccd1 vccd1 net1358 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_128_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout371 _06738_ vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__clkbuf_4
Xfanout1369 net1430 vssd1 vssd1 vccd1 vccd1 net1369 sky130_fd_sc_hd__buf_2
X_16740_ clknet_leaf_84_wb_clk_i _02427_ _00723_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout382 _03651_ vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__clkbuf_8
Xfanout393 net394 vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__clkbuf_8
X_13952_ _04220_ _04237_ _04239_ vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__and3_4
XFILLER_0_17_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10125__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12903_ net356 _03676_ _03677_ net869 net1663 vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__a32o_1
XANTENNA__10676__A1 _07015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16671_ clknet_leaf_41_wb_clk_i _02358_ _00654_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13883_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[9\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[7\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[6\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__or4b_1
XANTENNA__11904__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15622_ net1382 vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__inv_2
XANTENNA__09818__A0 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12834_ net2347 net188 net379 vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__mux2_1
XANTENNA__08338__X _04678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15553_ net1278 vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12765_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] net1060 net363 _03604_
+ vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__a22o_1
XANTENNA__09601__C net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10979__A2 _06590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14504_ net1353 vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__inv_2
X_11716_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] _07800_ vssd1 vssd1 vccd1
+ vccd1 _07910_ sky130_fd_sc_hd__nor2_1
X_15484_ net1246 vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__inv_2
X_12696_ net1950 net204 net383 vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17223_ clknet_leaf_105_wb_clk_i _02910_ _01206_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14435_ net1305 vssd1 vssd1 vccd1 vccd1 _00229_ sky130_fd_sc_hd__inv_2
XANTENNA__12735__S net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11647_ net1804 net203 net499 vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput13 DAT_I[1] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_840 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17154_ clknet_leaf_78_wb_clk_i _02841_ _01137_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput24 DAT_I[2] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
Xinput35 gpio_in[17] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_1
X_14366_ net1195 vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11578_ net575 _07793_ _07794_ vssd1 vssd1 vccd1 vccd1 _07795_ sky130_fd_sc_hd__and3_1
Xinput46 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08514__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput57 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_1
Xinput68 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__clkbuf_1
X_16105_ clknet_leaf_138_wb_clk_i _01880_ _00093_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[12\]
+ sky130_fd_sc_hd__dfrtp_4
X_13317_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[21\] net826 _03795_ _03797_
+ vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__o22a_1
Xhold808 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2343 sky130_fd_sc_hd__dlygate4sd3_1
X_17085_ clknet_leaf_64_wb_clk_i _02772_ _01068_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10529_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[31\] net674 net646 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[31\]
+ _06868_ vssd1 vssd1 vccd1 vccd1 _06869_ sky130_fd_sc_hd__a221o_1
Xhold819 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2354 sky130_fd_sc_hd__dlygate4sd3_1
X_14297_ net1329 vssd1 vssd1 vccd1 vccd1 _00091_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16036_ clknet_leaf_133_wb_clk_i _01830_ _00030_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09349__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13248_ net2521 net354 net350 team_01_WB.instance_to_wrap.cpu.f0.i\[2\] vssd1 vssd1
+ vccd1 vccd1 _01902_ sky130_fd_sc_hd__a22o_1
XANTENNA__09048__C net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12470__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13179_ net1549 net850 net842 vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__a21o_1
XANTENNA__14251__A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08887__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09345__A net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18006__1508 vssd1 vssd1 vccd1 vccd1 _18006__1508/HI net1508 sky130_fd_sc_hd__conb_1
Xhold1508 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net3043 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17987_ net1502 vssd1 vssd1 vccd1 vccd1 la_data_out[29] sky130_fd_sc_hd__buf_2
Xhold1519 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net3054 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_88_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16938_ clknet_leaf_33_wb_clk_i _02625_ _00921_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09521__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16869_ clknet_leaf_50_wb_clk_i _02556_ _00852_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11814__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09410_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[27\] net695 net662 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__a22o_1
XANTENNA__10938__B _07277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09341_ net598 _05678_ _05680_ vssd1 vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_62_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15810__A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09272_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[20\] net683 _05611_
+ net705 vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__a211o_1
XFILLER_0_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_115_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_115_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13369__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08223_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[58\] net2761 net1053 vssd1 vssd1
+ vccd1 vccd1 _03464_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12645__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout227_A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09588__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08154_ net1759 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[119\] net1048 vssd1 vssd1
+ vccd1 vccd1 _03533_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08085_ _04515_ _04523_ _04537_ _04557_ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__or4_1
XFILLER_0_141_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1136_A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12380__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1303_A net1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08987_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[8\] net661 _05325_ _05326_
+ net705 vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__a2111oi_1
XANTENNA_fanout763_A net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout384_X net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10107__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10658__A1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09512__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11009__B net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout930_A net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout649_X net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08720__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09608_ net996 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[24\] net982 vssd1
+ vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10880_ _05566_ _06708_ net368 vssd1 vssd1 vccd1 vccd1 _07220_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_51_Left_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09539_ net1152 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[28\] net969
+ vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__and3_1
XANTENNA__09276__A1 net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08079__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout816_X net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12550_ net2391 net309 net403 vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__mux2_1
XANTENNA__11083__B2 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11501_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[12\] _07756_ vssd1 vssd1 vccd1
+ vccd1 _07778_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12481_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[7\] net276 net412 vssd1
+ vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11312__X _07650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14220_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[12\] vssd1 vssd1 vccd1
+ vccd1 _02267_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11432_ team_01_WB.instance_to_wrap.cpu.f0.i\[6\] _07675_ net610 team_01_WB.instance_to_wrap.cpu.f0.i\[11\]
+ vssd1 vssd1 vccd1 vccd1 _07741_ sky130_fd_sc_hd__a31o_1
XANTENNA__09579__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14055__B _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14151_ net1632 net604 _04435_ net1185 vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__o211a_1
X_11363_ team_01_WB.instance_to_wrap.cpu.f0.i\[18\] team_01_WB.instance_to_wrap.cpu.f0.i\[17\]
+ _07690_ vssd1 vssd1 vccd1 vccd1 _07692_ sky130_fd_sc_hd__and3_1
X_13102_ net56 net55 net58 net57 vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__or4_1
X_10314_ net1129 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[18\] net951
+ vssd1 vssd1 vccd1 vccd1 _06654_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_60_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14082_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[76\] _04235_ _04268_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[76\]
+ vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11294_ _04714_ _07627_ _04734_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1
+ vssd1 vccd1 vccd1 _07634_ sky130_fd_sc_hd__a211o_1
X_17910_ net1521 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
X_13033_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[53\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[61\]
+ net859 vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__mux2_1
X_10245_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[9\] net777 net754 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06585_ sky130_fd_sc_hd__a22o_1
XANTENNA__12290__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1100 net1103 vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12886__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1111 net1113 vssd1 vssd1 vccd1 vccd1 net1111 sky130_fd_sc_hd__clkbuf_2
X_10176_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[10\] net780 _06514_
+ _06515_ vssd1 vssd1 vccd1 vccd1 _06516_ sky130_fd_sc_hd__a211o_1
XANTENNA__10897__A1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09751__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1122 net1123 vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__buf_2
X_17841_ clknet_leaf_121_wb_clk_i _03517_ _01781_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[111\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1133 net1134 vssd1 vssd1 vccd1 vccd1 net1133 sky130_fd_sc_hd__buf_2
Xfanout1144 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[19\] vssd1 vssd1 vccd1 vccd1
+ net1144 sky130_fd_sc_hd__buf_2
Xfanout1155 net1156 vssd1 vssd1 vccd1 vccd1 net1155 sky130_fd_sc_hd__buf_2
Xfanout1166 net1167 vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10104__A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14984_ net1374 vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__inv_2
X_17772_ clknet_leaf_92_wb_clk_i _03448_ _01712_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[42\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1177 net1178 vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__clkbuf_2
Xfanout1188 net1207 vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__buf_4
Xfanout190 net191 vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1199 net1200 vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10649__A1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13935_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[0\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__and2b_2
X_16723_ clknet_leaf_18_wb_clk_i _02410_ _00706_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_16654_ clknet_leaf_26_wb_clk_i _02341_ _00637_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13866_ net1178 net1065 net1709 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[27\]
+ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_83_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08509__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15605_ net1275 vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__inv_2
X_12817_ net1891 net641 net609 _03640_ vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__a22o_1
X_16585_ clknet_leaf_38_wb_clk_i _02272_ _00568_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[17\]
+ sky130_fd_sc_hd__dfrtp_4
X_13797_ _04175_ _04178_ vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15536_ net1272 vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__inv_2
X_12748_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] net1062 net365 _03592_
+ vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12810__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15467_ net1423 vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__inv_2
XANTENNA__12465__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12679_ net1929 net278 net388 vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08490__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17206_ clknet_leaf_30_wb_clk_i _02893_ _01189_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14418_ net1305 vssd1 vssd1 vccd1 vccd1 _00212_ sky130_fd_sc_hd__inv_2
X_15398_ net1400 vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17137_ clknet_leaf_113_wb_clk_i _02824_ _01120_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_14349_ net1333 vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold605 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2140 sky130_fd_sc_hd__dlygate4sd3_1
Xwire591 _04880_ vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__clkbuf_1
Xhold616 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2151 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold627 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2173 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold649 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2184 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17068_ clknet_leaf_16_wb_clk_i _02755_ _01051_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09990__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_51_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08910_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[2\] net671 _05229_ _05239_
+ _05246_ vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11809__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16019_ net1339 vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09890_ net1152 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[5\] net953 vssd1
+ vssd1 vccd1 vccd1 _06230_ sky130_fd_sc_hd__and3_1
XANTENNA__12877__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10888__A1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08841_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[1\] net694 _05156_ _05157_
+ _05170_ vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_85_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09506__C net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1305 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[78\] vssd1 vssd1 vccd1 vccd1
+ net2840 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11892__X _07949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1316 _02150_ vssd1 vssd1 vccd1 vccd1 net2851 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1327 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2862 sky130_fd_sc_hd__dlygate4sd3_1
X_08772_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[11\] net729 _05111_ net1080 vssd1
+ vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__a22o_1
Xhold1338 _03516_ vssd1 vssd1 vccd1 vccd1 net2873 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1349 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2884 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_108_Left_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_144_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08702__B1 _05041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout344_A _04748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1086_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09324_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[24\] net686 net673 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10812__A1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09255_ net598 _05591_ _05593_ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__o21a_1
XFILLER_0_63_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12375__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout511_A _05963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout609_A _03583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_90_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08206_ net2565 net2418 net1054 vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_117_Left_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11499__B _07756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09186_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[16\] net684 _05523_
+ _05524_ _05525_ vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12565__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08137_ _04467_ team_01_WB.instance_to_wrap.cpu.f0.num\[28\] team_01_WB.instance_to_wrap.cpu.f0.num\[21\]
+ _04473_ _04596_ vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__a221o_1
XANTENNA__13995__A _04152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10576__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1041_X net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07993__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_83_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09981__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08068_ _04514_ _04532_ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout880_A net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11719__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout599_X net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_12_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_105_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12868__A2 _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10030_ net994 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[0\] net981 vssd1
+ vssd1 vccd1 vccd1 _06370_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09733__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout766_X net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_126_Left_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11981_ net2474 net252 net474 vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout933_X net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13720_ _04107_ _04129_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[11\]
+ sky130_fd_sc_hd__nor2_1
X_10932_ _05338_ _06563_ vssd1 vssd1 vccd1 vccd1 _07272_ sky130_fd_sc_hd__or2_1
XANTENNA__08329__A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13651_ _03877_ _03879_ vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__xnor2_1
X_10863_ _06980_ _07132_ _07202_ _06920_ vssd1 vssd1 vccd1 vccd1 _07203_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_155_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12602_ net2349 net233 net395 vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16370_ clknet_leaf_101_wb_clk_i _02124_ _00353_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[93\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__13889__B _04146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13582_ net721 _07541_ net1074 vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__o21a_1
XFILLER_0_66_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10794_ _06963_ _07122_ _07133_ _07054_ _07131_ vssd1 vssd1 vccd1 vccd1 _07134_ sky130_fd_sc_hd__a221o_1
XFILLER_0_109_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08990__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15321_ net1233 vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__inv_2
X_12533_ net2727 net244 net404 vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_135_Left_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12285__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15252_ net1378 vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__inv_2
X_12464_ net2658 net272 net413 vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16054__Q team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14203_ net2384 vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__clkbuf_1
X_11415_ team_01_WB.instance_to_wrap.cpu.f0.i\[18\] _07705_ vssd1 vssd1 vccd1 vccd1
+ _07731_ sky130_fd_sc_hd__or2_1
XANTENNA__11202__B _07520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15183_ net1296 vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_750 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10567__A0 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12395_ net2339 net210 net419 vssd1 vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__mux2_1
XANTENNA__08999__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14134_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[31\] _04243_ _04261_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[119\]
+ _04418_ vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__a221o_1
X_11346_ team_01_WB.instance_to_wrap.cpu.f0.i\[5\] team_01_WB.instance_to_wrap.cpu.f0.i\[4\]
+ _07674_ vssd1 vssd1 vccd1 vccd1 _07675_ sky130_fd_sc_hd__and3_1
XANTENNA__09972__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14065_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[19\] _04259_ _04349_ _04351_
+ _04353_ vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__a2111o_1
X_11277_ _05595_ net331 _07354_ net336 net369 vssd1 vssd1 vccd1 vccd1 _07617_ sky130_fd_sc_hd__a221o_1
XANTENNA__10319__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13016_ net2949 net2912 net854 vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10228_ _06566_ _06567_ vssd1 vssd1 vccd1 vccd1 _06568_ sky130_fd_sc_hd__nand2_1
XANTENNA__09724__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_135_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17824_ clknet_leaf_120_wb_clk_i net2731 _01764_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[94\]
+ sky130_fd_sc_hd__dfrtp_1
X_10159_ _06497_ _06498_ net340 vssd1 vssd1 vccd1 vccd1 _06499_ sky130_fd_sc_hd__a21oi_1
Xhold2 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[7\] vssd1 vssd1 vccd1 vccd1 net1537
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17755_ clknet_leaf_92_wb_clk_i net2430 _01695_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_14967_ net1243 vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__inv_2
X_16706_ clknet_leaf_78_wb_clk_i _02393_ _00689_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10098__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13918_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[12\] _04212_ net571 vssd1
+ vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_18_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14898_ net1290 vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__inv_2
X_17686_ clknet_leaf_128_wb_clk_i _03370_ _01627_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09910__X _06250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09061__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16637_ clknet_leaf_69_wb_clk_i _02324_ _00620_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13849_ net1179 net1066 net3188 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[10\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16568_ clknet_leaf_27_wb_clk_i _02255_ _00551_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_71_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12795__A1 _07207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13992__B1 _04266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15519_ net1314 vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__inv_2
XANTENNA__12195__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16499_ clknet_leaf_156_wb_clk_i _02253_ _00482_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09040_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] _04846_ net593 vssd1 vssd1
+ vccd1 vccd1 _05380_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_72_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold402 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1937 sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1948 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10022__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold424 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1959 sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1970 sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[120\] vssd1 vssd1 vccd1 vccd1
+ net1981 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13441__A_N _05456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold457 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1992 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold468 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2003 sky130_fd_sc_hd__dlygate4sd3_1
X_09942_ net377 _05264_ vssd1 vssd1 vccd1 vccd1 _06282_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_74_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold479 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2014 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout904 _04785_ vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_74_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout915 net916 vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout926 net928 vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__buf_2
XANTENNA__09715__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09873_ _06198_ _06210_ _06211_ _06212_ vssd1 vssd1 vccd1 vccd1 _06213_ sky130_fd_sc_hd__or4_1
Xfanout937 net938 vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__clkbuf_2
Xfanout948 net950 vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__buf_4
XANTENNA_fanout294_A net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout959 net961 vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__buf_4
X_08824_ net1105 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[1\] net889 vssd1
+ vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_5_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1102 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[32\] vssd1 vssd1 vccd1 vccd1
+ net2637 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1113 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2648 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1124 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2659 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1001_A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1135 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2670 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2681 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09533__A net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08755_ net1099 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[4\] net924 vssd1
+ vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__and3_1
Xhold1157 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2692 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout461_A _07955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1168 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1179 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[31\] vssd1 vssd1 vccd1 vccd1
+ net2714 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout559_A net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10089__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08686_ net1006 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[7\] net882 vssd1
+ vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_130_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_130_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_120_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout726_A net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout347_X net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1089_X net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08436__X _04776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12786__A1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09307_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[22\] net674 _05621_
+ _05631_ _05639_ vssd1 vssd1 vccd1 vccd1 _05647_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13983__B1 _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10618__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09238_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[21\] net696 net694 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[21\]
+ _05577_ vssd1 vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08315__C net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11022__B net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09169_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[16\] net652 _05506_
+ _05507_ _05508_ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10549__A0 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09403__A1 net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11200_ _06963_ _07054_ _07324_ net557 vssd1 vssd1 vccd1 vccd1 _07540_ sky130_fd_sc_hd__o22a_1
XANTENNA__11210__A1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09708__A net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10013__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12180_ net2443 net280 net448 vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout883_X net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11131_ _06399_ _06401_ vssd1 vssd1 vccd1 vccd1 _07471_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold980 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2515 sky130_fd_sc_hd__dlygate4sd3_1
Xhold991 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2526 sky130_fd_sc_hd__dlygate4sd3_1
X_11062_ _07394_ _07398_ _07400_ _07401_ vssd1 vssd1 vccd1 vccd1 _07402_ sky130_fd_sc_hd__a211o_1
X_10013_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[1\] net780 net761 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06353_ sky130_fd_sc_hd__a22o_1
X_15870_ net1203 vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__inv_2
XANTENNA__08985__C net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14821_ net1262 vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__inv_2
XANTENNA_input22_A DAT_I[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09443__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10589__A net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17540_ clknet_leaf_73_wb_clk_i _03227_ _01523_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_14752_ net1187 vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__inv_2
XANTENNA__11277__B2 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11964_ net2632 net211 net471 vssd1 vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__mux2_1
X_13703_ _04104_ _04119_ _04122_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[7\]
+ sky130_fd_sc_hd__and3_1
X_17471_ clknet_leaf_45_wb_clk_i _03158_ _01454_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10915_ net374 net373 net371 _06158_ net539 net546 vssd1 vssd1 vccd1 vccd1 _07255_
+ sky130_fd_sc_hd__mux4_1
X_14683_ net1306 vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__inv_2
XANTENNA__08693__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11895_ net2395 _07831_ net481 vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11912__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15180__A net1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_143_Left_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16422_ clknet_leaf_135_wb_clk_i _02176_ _00405_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13634_ net722 _07290_ net1073 vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__o21a_1
X_10846_ net528 _06921_ _06972_ _06978_ _07185_ vssd1 vssd1 vccd1 vccd1 _07186_ sky130_fd_sc_hd__o311ai_2
X_16353_ clknet_leaf_118_wb_clk_i _02107_ _00336_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[76\]
+ sky130_fd_sc_hd__dfstp_1
X_13565_ net720 _07135_ net1073 vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__o21a_1
XANTENNA__13412__B _05224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10777_ net509 net508 net507 net505 net549 net542 vssd1 vssd1 vccd1 vccd1 _07117_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_27_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15304_ net1375 vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__inv_2
X_12516_ net1751 net294 net410 vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__mux2_1
XANTENNA__10252__A2 _05338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16284_ clknet_leaf_124_wb_clk_i _02038_ _00267_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13496_ net185 _03955_ _03956_ net723 vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__a211o_1
X_15235_ net1251 vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__inv_2
X_12447_ net2826 net302 net416 vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15166_ net1316 vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__inv_2
X_12378_ net2399 net225 net423 vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14117_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[110\] _04264_ _04400_ _04402_
+ vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__a211o_1
X_11329_ _04547_ _07653_ _07662_ net1176 vssd1 vssd1 vccd1 vccd1 _07663_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15097_ net1237 vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_52_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10490__C net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14048_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[67\] _04233_ _04260_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[59\]
+ vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__a22o_1
XANTENNA__09056__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11504__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12701__A1 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15355__A net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08895__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17807_ clknet_leaf_100_wb_clk_i _03483_ _01747_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[77\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_141_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15999_ net1413 vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08540_ _04871_ _04872_ _04878_ _04879_ vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__nor4_1
XANTENNA__11268__B2 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17738_ clknet_leaf_123_wb_clk_i _03414_ _01678_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09330__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08471_ net1109 net880 vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17669_ clknet_leaf_157_wb_clk_i _03354_ _01610_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11822__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12768__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09023_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[9\] net688 _05342_ _05347_
+ _05362_ vssd1 vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_142_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12653__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout307_A _07935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09397__B1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1049_A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold210 team_01_WB.instance_to_wrap.a1.ADR_I\[27\] vssd1 vssd1 vccd1 vccd1 net1745
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09936__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold221 net150 vssd1 vssd1 vccd1 vccd1 net1756 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08432__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold232 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1767 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold243 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1778 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12940__A1 _05005_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold254 _02154_ vssd1 vssd1 vccd1 vccd1 net1789 sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[121\] vssd1 vssd1 vccd1 vccd1
+ net1800 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 _03341_ vssd1 vssd1 vccd1 vccd1 net1811 sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1822 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1216_A net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout701 _04758_ vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__buf_8
Xhold298 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1833 sky130_fd_sc_hd__dlygate4sd3_1
X_09925_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[4\] net792 _06262_ _06263_
+ _06264_ vssd1 vssd1 vccd1 vccd1 _06265_ sky130_fd_sc_hd__a2111o_1
XANTENNA__14142__B1 _04265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout723 net728 vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__clkbuf_4
Xfanout734 net736 vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__clkbuf_8
Xfanout745 net748 vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout676_A _04790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout756 _04675_ vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__clkbuf_4
X_09856_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[12\] net796 net778 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06196_ sky130_fd_sc_hd__a22o_1
Xfanout767 _04673_ vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__clkbuf_4
Xfanout778 _04666_ vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1004_X net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout789 net790 vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__clkbuf_8
X_08807_ net1093 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[0\] net879 vssd1
+ vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__and3_1
Xclkbuf_4_8__f_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_8__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_09787_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[15\] net765 vssd1 vssd1
+ vccd1 vccd1 _06127_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout464_X net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout843_A net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08738_ net1099 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[4\] net884 vssd1
+ vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13653__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09321__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08669_ net1006 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[7\] net896 vssd1
+ vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout631_X net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10700_ net535 _06955_ vssd1 vssd1 vccd1 vccd1 _07040_ sky130_fd_sc_hd__or2_1
X_11680_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[15\] net713 vssd1 vssd1 vccd1
+ vccd1 _07881_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12759__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10631_ net514 _06857_ vssd1 vssd1 vccd1 vccd1 _06971_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08326__B net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10234__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13350_ team_01_WB.instance_to_wrap.cpu.f0.i\[11\] _07677_ vssd1 vssd1 vccd1 vccd1
+ _03823_ sky130_fd_sc_hd__or2_1
X_10562_ _06900_ _06901_ vssd1 vssd1 vccd1 vccd1 _06902_ sky130_fd_sc_hd__or2_2
X_12301_ net2733 net200 net432 vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13281_ _07650_ _03767_ _03769_ net825 net3155 vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__o32a_1
XANTENNA__12563__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10493_ net1130 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[31\] net965 vssd1
+ vssd1 vccd1 vccd1 _06833_ sky130_fd_sc_hd__and3b_1
X_15020_ net1257 vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__inv_2
X_12232_ net3030 net207 net441 vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__mux2_1
XANTENNA__12931__A1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12163_ net2755 net245 net449 vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__mux2_1
XANTENNA__10942__A0 _06636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09725__X _06065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11114_ _07452_ _07453_ net540 vssd1 vssd1 vccd1 vccd1 _07454_ sky130_fd_sc_hd__mux2_1
XANTENNA__14133__B1 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16971_ clknet_leaf_8_wb_clk_i _02658_ _00954_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_12094_ net3138 net220 net457 vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__mux2_1
XANTENNA__11907__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11045_ net541 _07011_ _06366_ vssd1 vssd1 vccd1 vccd1 _07385_ sky130_fd_sc_hd__o21ai_1
X_15922_ net1353 vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09173__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15853_ net1334 vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__inv_2
XANTENNA__09604__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14804_ net1379 vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12996_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[90\] net2898 net863 vssd1 vssd1
+ vccd1 vccd1 _02129_ sky130_fd_sc_hd__mux2_1
X_15784_ net1203 vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17523_ clknet_leaf_18_wb_clk_i _03210_ _01506_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11947_ net2179 net251 net478 vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14735_ net1198 vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12738__S net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11642__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14666_ net1305 vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__inv_2
XANTENNA__11670__A1 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17454_ clknet_leaf_28_wb_clk_i _03141_ _01437_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11878_ net2392 net256 net484 vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__mux2_1
XANTENNA__08517__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13617_ net721 _07207_ net1075 vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__o21a_1
X_16405_ clknet_leaf_124_wb_clk_i _02159_ _00388_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10829_ _07064_ _07099_ _07167_ _07168_ vssd1 vssd1 vccd1 vccd1 _07169_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_45_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17385_ clknet_leaf_38_wb_clk_i _03072_ _01368_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14597_ net1362 vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13548_ net720 _07154_ net1073 vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__o21a_1
X_16336_ clknet_leaf_95_wb_clk_i net2481 _00319_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16267_ clknet_leaf_141_wb_clk_i net1599 _00255_ vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13479_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] _05679_ vssd1 vssd1
+ vccd1 vccd1 _03940_ sky130_fd_sc_hd__xor2_1
XANTENNA__10782__A net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12473__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14254__A net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13175__A1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18006_ net1508 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__buf_2
X_15218_ net1267 vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__inv_2
XANTENNA__09379__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09918__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16198_ clknet_leaf_159_wb_clk_i _01958_ _00186_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_93_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15149_ net1265 vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10933__A0 _06919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14124__B1 _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07971_ team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1 _04469_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_10_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11817__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09710_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[21\] net795 _06038_ _06039_
+ _06040_ vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10721__S net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09083__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09641_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[23\] net811 net742 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15813__A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09572_ net1149 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[25\] net976
+ vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_69_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08523_ net1079 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[18\] net906
+ vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__and3_1
XANTENNA__12648__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08657__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11110__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13650__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08454_ net1021 net898 vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__and2_1
XANTENNA__10464__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08385_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout424_A net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_154_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12383__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09006_ net1012 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[9\] net900 vssd1
+ vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__and3_1
XANTENNA__09909__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1121_X net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09790__B1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14115__B1 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout520 _05260_ vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout679_X net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout531 net532 vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__buf_2
Xfanout542 _05189_ vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__buf_2
X_09908_ net770 _06240_ _06244_ _06247_ vssd1 vssd1 vccd1 vccd1 _06248_ sky130_fd_sc_hd__or4_2
Xfanout553 net554 vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__buf_2
Xfanout564 net566 vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__buf_2
Xfanout575 _07792_ vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__buf_2
Xfanout586 net587 vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__buf_2
X_09839_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[13\] net815 net738 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06179_ sky130_fd_sc_hd__a22o_1
Xfanout597 net599 vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__clkbuf_8
X_12850_ net2927 net229 net380 vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__mux2_1
X_17959__1474 vssd1 vssd1 vccd1 vccd1 _17959__1474/HI net1474 sky130_fd_sc_hd__conb_1
X_11801_ net2189 net202 net491 vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__mux2_1
X_12781_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] net1062 net364 _03615_
+ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__a22o_1
Xclkbuf_3_1_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12558__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14520_ net1352 vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__inv_2
X_11732_ net715 _07507_ net612 vssd1 vssd1 vccd1 vccd1 _07923_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10455__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08337__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14451_ net1227 vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11663_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] _07812_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\]
+ vssd1 vssd1 vccd1 vccd1 _07868_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_153_Right_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13402_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\]
+ net596 vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__and3_1
XFILLER_0_153_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10207__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10614_ net546 _06366_ vssd1 vssd1 vccd1 vccd1 _06954_ sky130_fd_sc_hd__nor2_1
X_17170_ clknet_leaf_144_wb_clk_i _02857_ _01153_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_14382_ net1193 vssd1 vssd1 vccd1 vccd1 _00176_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09073__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11594_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] _07809_ vssd1 vssd1
+ vccd1 vccd1 _07811_ sky130_fd_sc_hd__nand2_1
Xwire921 _04775_ vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16121_ clknet_leaf_136_wb_clk_i _01896_ _00109_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[28\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_52_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13333_ team_01_WB.instance_to_wrap.cpu.f0.i\[15\] _07682_ net826 vssd1 vssd1 vccd1
+ vccd1 _03810_ sky130_fd_sc_hd__o21a_1
X_10545_ _06883_ _06884_ vssd1 vssd1 vccd1 vccd1 _06885_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12293__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08820__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap709 _04729_ vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__buf_1
XFILLER_0_51_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09168__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16052_ clknet_leaf_15_wb_clk_i _01845_ _00040_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13264_ net587 _03750_ _03755_ net564 _04466_ vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__a221oi_1
X_10476_ net512 _05933_ net511 _05964_ vssd1 vssd1 vccd1 vccd1 _06816_ sky130_fd_sc_hd__a22o_1
XANTENNA__08072__A team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_121_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15003_ net1254 vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__inv_2
XANTENNA__12904__A1 _05591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11707__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12215_ net2016 net276 net444 vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13195_ net14 net835 net628 net2608 vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__o22a_1
XANTENNA__10915__A0 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14106__B1 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12146_ net3156 net252 net454 vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__mux2_1
XANTENNA__09781__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11637__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16954_ clknet_leaf_78_wb_clk_i _02641_ _00937_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12077_ net2353 net255 net460 vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__mux2_1
X_11028_ _07366_ _07367_ vssd1 vssd1 vccd1 vccd1 _07368_ sky130_fd_sc_hd__and2_1
X_15905_ net1402 vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__inv_2
X_16885_ clknet_leaf_118_wb_clk_i _02572_ _00868_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15836_ net1330 vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15767_ net1199 vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__inv_2
XANTENNA__17621__Q team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12468__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12979_ net2532 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[115\] net862 vssd1 vssd1
+ vccd1 vccd1 _02146_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17506_ clknet_leaf_56_wb_clk_i _03193_ _01489_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_14718_ net1186 vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__inv_2
XANTENNA__11643__A1 _07111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15698_ net1289 vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17437_ clknet_leaf_69_wb_clk_i _03124_ _01420_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_145_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14649_ net1249 vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_16 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_28_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_27 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_38 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08170_ net3005 net2824 net1047 vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__mux2_1
X_17368_ clknet_leaf_61_wb_clk_i _03055_ _01351_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_49 _03654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16319_ clknet_leaf_91_wb_clk_i net2047 _00302_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08811__A2 _05150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17299_ clknet_leaf_24_wb_clk_i _02986_ _01282_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_132_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__buf_2
XANTENNA__09509__C net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__buf_2
XFILLER_0_88_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput123 net123 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__buf_2
XFILLER_0_140_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15808__A net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput134 net134 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__buf_2
Xoutput145 net145 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__buf_2
XANTENNA__13182__A_N net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput156 net156 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
XANTENNA__09365__X _05705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput167 net167 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__clkbuf_4
XANTENNA__09772__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput178 net178 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__clkbuf_4
XANTENNA__08710__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10382__A1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout374_A _06129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09624_ _05682_ _05734_ vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_108_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09541__A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13084__A0 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09555_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[28\] net792 net768 _05883_
+ _05894_ vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__a2111o_1
Xclkbuf_leaf_37_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12378__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout541_A net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout639_A _03572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13623__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08506_ net711 _04838_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__or2_2
XANTENNA__11634__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09486_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[30\] net676 net648 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_156_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08437_ net1004 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[23\] net917 vssd1
+ vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_22_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_156_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout427_X net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1169_X net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08368_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[2\] _04623_ _04626_ vssd1 vssd1
+ vccd1 vccd1 _04708_ sky130_fd_sc_hd__nor3_2
XFILLER_0_34_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08299_ net991 net975 vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10330_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[18\] net763 net622 vssd1
+ vssd1 vccd1 vccd1 _06670_ sky130_fd_sc_hd__o21a_1
XFILLER_0_132_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout796_X net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11030__B net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10261_ net339 _06593_ _06566_ vssd1 vssd1 vccd1 vccd1 _06601_ sky130_fd_sc_hd__a21boi_2
XANTENNA__12841__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12000_ net2378 net272 net468 vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__mux2_1
XANTENNA__09275__X _05615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10192_ _06530_ _06531_ vssd1 vssd1 vccd1 vccd1 _06532_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout963_X net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1304 net38 vssd1 vssd1 vccd1 vccd1 net1304 sky130_fd_sc_hd__buf_4
Xfanout1315 net1322 vssd1 vssd1 vccd1 vccd1 net1315 sky130_fd_sc_hd__clkbuf_4
Xfanout1326 net1327 vssd1 vssd1 vccd1 vccd1 net1326 sky130_fd_sc_hd__clkbuf_4
Xfanout1337 net1344 vssd1 vssd1 vccd1 vccd1 net1337 sky130_fd_sc_hd__buf_2
Xfanout350 _03742_ vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__buf_2
Xfanout1348 net1349 vssd1 vssd1 vccd1 vccd1 net1348 sky130_fd_sc_hd__buf_4
Xfanout361 _03653_ vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__buf_4
Xfanout1359 net1362 vssd1 vssd1 vccd1 vccd1 net1359 sky130_fd_sc_hd__buf_2
Xfanout372 _06465_ vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__buf_2
X_13951_ _04225_ _04242_ vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__nor2_4
Xfanout383 _03570_ vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__buf_6
XANTENNA__08869__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10125__B2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout394 _03568_ vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__buf_6
X_12902_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[22\] net1037 vssd1 vssd1 vccd1
+ vccd1 _03677_ sky130_fd_sc_hd__or2_1
X_16670_ clknet_leaf_80_wb_clk_i _02357_ _00653_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13882_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[4\]
+ _04188_ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__and3_1
XANTENNA__08993__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15621_ net1289 vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__inv_2
X_12833_ net576 _07794_ _07945_ vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__and3_1
XANTENNA__12288__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09818__A1 _06157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10428__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12764_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[21\] _07621_ net1034 vssd1 vssd1
+ vccd1 vccd1 _03604_ sky130_fd_sc_hd__mux2_1
X_15552_ net1239 vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16057__Q team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10979__A3 _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11715_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[8\] _07290_ net714 vssd1 vssd1
+ vccd1 vccd1 _07909_ sky130_fd_sc_hd__mux2_1
X_14503_ net1400 vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__inv_2
X_15483_ net1248 vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__inv_2
X_12695_ net2613 net275 net385 vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__mux2_1
XANTENNA__11920__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17222_ clknet_leaf_72_wb_clk_i _02909_ _01205_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11646_ _07852_ _07854_ net611 vssd1 vssd1 vccd1 vccd1 _07855_ sky130_fd_sc_hd__mux2_4
X_14434_ net1307 vssd1 vssd1 vccd1 vccd1 _00228_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput14 DAT_I[20] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
X_17153_ clknet_leaf_55_wb_clk_i _02840_ _01136_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput25 DAT_I[30] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
X_14365_ net1206 vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput36 gpio_in[18] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_1
X_11577_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\] team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\]
+ vssd1 vssd1 vccd1 vccd1 _07794_ sky130_fd_sc_hd__and2_2
XFILLER_0_80_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput47 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_1
X_13316_ net564 _07708_ _03796_ net828 vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__a31o_1
Xinput58 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_1
X_16104_ clknet_leaf_127_wb_clk_i _01879_ _00092_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_17084_ clknet_leaf_58_wb_clk_i _02771_ _01067_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput69 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__dlymetal6s2s_1
X_10528_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[31\] net683 net667 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06868_ sky130_fd_sc_hd__a22o_1
Xhold809 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2344 sky130_fd_sc_hd__dlygate4sd3_1
X_14296_ net1329 vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__inv_2
XFILLER_0_149_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_41_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13247_ net2579 net353 net349 team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1
+ vccd1 vccd1 _01903_ sky130_fd_sc_hd__a22o_1
X_16035_ clknet_leaf_136_wb_clk_i _01829_ _00029_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10459_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[26\] net812 net775 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06799_ sky130_fd_sc_hd__a22o_1
XANTENNA__13550__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09754__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09626__A net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13178_ net3152 net847 net634 vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__a21o_1
X_12129_ net2174 net210 net451 vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17986_ net1501 vssd1 vssd1 vccd1 vccd1 la_data_out[28] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_36_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1509 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net3044 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13302__A1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16937_ clknet_leaf_35_wb_clk_i _02624_ _00920_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09064__C net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11864__A1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16868_ clknet_leaf_73_wb_clk_i _02555_ _00851_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_15819_ net1190 vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12198__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16799_ clknet_leaf_43_wb_clk_i _02486_ _00782_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_09340_ net600 _05679_ vssd1 vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__or2_2
XANTENNA__11616__A1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10300__A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12813__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09271_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[20\] net662 net658 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_16_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10794__X _07134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11830__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08222_ net2661 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[51\] net1054 vssd1 vssd1
+ vccd1 vccd1 _03465_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_80_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_28_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08705__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14030__A2 _04230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08153_ team_01_WB.instance_to_wrap.cpu.f0.read_i net827 _00020_ vssd1 vssd1 vccd1
+ vccd1 _03534_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_151_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_155_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_155_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_71_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08084_ _04528_ _04532_ _04527_ vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12661__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17958__1473 vssd1 vssd1 vccd1 vccd1 _17958__1473/HI net1473 sky130_fd_sc_hd__conb_1
XFILLER_0_140_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1129_A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08440__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11552__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout491_A _07944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08986_ net1007 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[8\] net879 vssd1
+ vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__and3_1
XANTENNA__14097__A2 _04254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout756_A _04675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout377_X net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08439__X _04779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09607_ net996 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[24\] net949 vssd1
+ vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_123_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout923_A _04770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09702__C net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12804__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09538_ net1152 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[28\] net949
+ vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09276__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11025__B net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11083__A2 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout711_X net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09469_ net1083 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[30\] net878
+ vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12836__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout809_X net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11500_ net1962 net876 _07758_ _07777_ vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__o22a_1
XFILLER_0_109_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12480_ net3129 net302 net412 vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09028__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14021__A2 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11431_ _07680_ _07701_ _07740_ net324 vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__o211a_1
XANTENNA__08334__B net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10043__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14150_ _04422_ _04431_ _04433_ _04434_ vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__or4_1
XANTENNA__14055__C _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11362_ team_01_WB.instance_to_wrap.cpu.f0.i\[17\] _07690_ vssd1 vssd1 vccd1 vccd1
+ _07691_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13101_ net47 net49 net48 net46 vssd1 vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__or4b_1
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10313_ _06650_ _06651_ _06652_ vssd1 vssd1 vccd1 vccd1 _06653_ sky130_fd_sc_hd__or3_1
XANTENNA__12571__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14081_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[124\] _04263_ _04264_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[108\]
+ _04368_ vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11293_ _07627_ _07629_ _07632_ vssd1 vssd1 vccd1 vccd1 _07633_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_131_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13032_ net2629 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[62\] net854 vssd1 vssd1
+ vccd1 vccd1 _02093_ sky130_fd_sc_hd__mux2_1
X_10244_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[9\] net823 net788 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06584_ sky130_fd_sc_hd__a22o_1
XANTENNA__08988__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11695__B net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input52_A wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09446__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11543__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1101 net1102 vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__clkbuf_2
Xfanout1112 net1113 vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__buf_1
XANTENNA_clkbuf_leaf_125_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17840_ clknet_leaf_120_wb_clk_i net2873 _01780_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[110\]
+ sky130_fd_sc_hd__dfrtp_1
X_10175_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[10\] _04659_ net738
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[10\] vssd1 vssd1 vccd1 vccd1
+ _06515_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1123 net1124 vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__buf_1
Xfanout1134 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[19\] vssd1 vssd1 vccd1 vccd1
+ net1134 sky130_fd_sc_hd__buf_2
XANTENNA__14088__A2 _04375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1145 net1151 vssd1 vssd1 vccd1 vccd1 net1145 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1156 net1157 vssd1 vssd1 vccd1 vccd1 net1156 sky130_fd_sc_hd__clkbuf_4
X_17771_ clknet_leaf_93_wb_clk_i _03447_ _01711_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[41\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1167 net1168 vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__buf_1
X_14983_ net1387 vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__inv_2
Xfanout1178 net1181 vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__buf_2
XANTENNA__11915__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1189 net1192 vssd1 vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__buf_4
Xfanout191 _07823_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__clkbuf_2
X_16722_ clknet_leaf_113_wb_clk_i _02409_ _00705_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13934_ _04224_ _04225_ vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__nor2_4
XFILLER_0_117_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09181__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16653_ clknet_leaf_68_wb_clk_i _02340_ _00636_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13865_ net1178 net1064 net2115 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[26\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_92_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15604_ net1378 vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__inv_2
X_12816_ net364 _03638_ _03639_ net1063 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__a32o_1
X_16584_ clknet_leaf_62_wb_clk_i _02271_ _00567_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13796_ _04177_ _04174_ _01836_ vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09267__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15535_ net1299 vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__inv_2
X_12747_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[26\] _07588_ net1036 vssd1 vssd1
+ vccd1 vccd1 _03592_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11650__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10282__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12678_ net2148 net301 net388 vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__mux2_1
X_15466_ net1284 vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__inv_2
XANTENNA__14012__A2 _04241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08525__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17205_ clknet_leaf_113_wb_clk_i _02892_ _01188_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11629_ _07819_ _07840_ vssd1 vssd1 vccd1 vccd1 _07841_ sky130_fd_sc_hd__nor2_1
X_14417_ net1323 vssd1 vssd1 vccd1 vccd1 _00211_ sky130_fd_sc_hd__inv_2
X_15397_ net1287 vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__inv_2
XANTENNA__10493__C net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09908__X _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17136_ clknet_leaf_146_wb_clk_i _02823_ _01119_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14348_ net1326 vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__inv_2
Xhold606 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2141 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09059__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10585__A1 _06882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwire581 _06705_ vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__clkbuf_2
Xhold617 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2152 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwire592 _04877_ vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__clkbuf_1
Xhold628 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2163 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12481__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14279_ net1336 vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_38_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17067_ clknet_leaf_9_wb_clk_i _02754_ _01050_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold639 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2174 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13523__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08898__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16018_ net1329 vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[1\] net663 _05159_ _05173_
+ _05174_ vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_55_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10888__A2 _07227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14079__A2 _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1306 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[94\] vssd1 vssd1 vccd1 vccd1
+ net2841 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08771_ _04708_ net725 net718 _04838_ vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__or4_2
Xhold1317 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2852 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17969_ net1484 vssd1 vssd1 vccd1 vccd1 la_data_out[11] sky130_fd_sc_hd__buf_2
Xhold1328 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2863 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1339 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2874 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_144_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08702__A1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10030__A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09258__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09323_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[24\] _04766_ net677
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[24\] vssd1 vssd1 vccd1 vccd1
+ _05663_ sky130_fd_sc_hd__a22o_1
XANTENNA__12656__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09254_ net597 _05591_ _05593_ vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_29_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1079_A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14003__A2 _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08205_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[76\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[68\]
+ net1045 vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09185_ net1091 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[16\] net917
+ vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_32_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout504_A _06779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1246_A net1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08136_ team_01_WB.instance_to_wrap.cpu.f0.i\[28\] _04494_ team_01_WB.instance_to_wrap.cpu.f0.num\[0\]
+ _04489_ _04605_ vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__a221o_1
XANTENNA__09818__X _06158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10576__A1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09430__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08067_ _04528_ _04539_ vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__nor2_1
XANTENNA__12391__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14172__A net1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1034_X net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13514__A1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_15__f_wb_clk_i_X clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout494_X net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_52_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout661_X net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08969_ net1088 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[8\] net888 vssd1
+ vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_125_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout759_X net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11980_ net2527 net226 net471 vssd1 vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__mux2_1
X_10931_ _05338_ _06563_ vssd1 vssd1 vccd1 vccd1 _07271_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout926_X net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08329__B net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10862_ net503 _07105_ net375 vssd1 vssd1 vccd1 vccd1 _07202_ sky130_fd_sc_hd__mux2_1
X_13650_ net988 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] _04083_ _04084_
+ vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__a22o_1
XANTENNA__09249__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12601_ net2993 net237 net395 vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13581_ net187 _04025_ _04026_ net727 vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__a211o_1
XFILLER_0_13_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10793_ net528 _07132_ _07119_ vssd1 vssd1 vccd1 vccd1 _07133_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13863__A_N net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12566__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12532_ net2134 net202 net403 vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__mux2_1
X_15320_ net1215 vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10594__B _06902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15251_ net1383 vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__inv_2
X_12463_ net2781 net207 net413 vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__mux2_1
XANTENNA__13202__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10016__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11414_ team_01_WB.instance_to_wrap.cpu.f0.i\[18\] _07691_ vssd1 vssd1 vccd1 vccd1
+ _07730_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14202_ net3012 vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15182_ net1300 vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__inv_2
XANTENNA__11202__C _07531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12394_ net2805 net214 net419 vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__mux2_1
XANTENNA__10567__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09421__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14133_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[47\] _04246_ _04252_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[111\]
+ vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11345_ team_01_WB.instance_to_wrap.cpu.f0.i\[3\] _07673_ vssd1 vssd1 vccd1 vccd1
+ _07674_ sky130_fd_sc_hd__and2_1
XFILLER_0_61_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09709__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09176__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14064_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[11\] _04253_ _04261_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[115\]
+ _04352_ vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__a221o_1
X_11276_ _06919_ _07354_ vssd1 vssd1 vccd1 vccd1 _07616_ sky130_fd_sc_hd__nor2_1
XANTENNA__09607__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16070__Q team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13015_ net2678 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[79\] net856 vssd1 vssd1
+ vccd1 vccd1 _02110_ sky130_fd_sc_hd__mux2_1
XANTENNA__08511__C net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10227_ _06562_ _06565_ vssd1 vssd1 vccd1 vccd1 _06567_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_33_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09463__X _05803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17823_ clknet_leaf_100_wb_clk_i _03499_ _01763_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[93\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10158_ net377 _05379_ net376 vssd1 vssd1 vccd1 vccd1 _06498_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_7_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[4\] vssd1 vssd1 vccd1 vccd1 net1538
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_50_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17754_ clknet_leaf_123_wb_clk_i _03430_ _01694_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10089_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[7\] net786 net782 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06429_ sky130_fd_sc_hd__a22o_1
X_14966_ net1256 vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_50_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16705_ clknet_leaf_55_wb_clk_i _02392_ _00688_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13917_ _04212_ net571 _04211_ vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_18_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17685_ clknet_leaf_128_wb_clk_i _03369_ _01626_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_14897_ net1423 vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_18_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16636_ clknet_leaf_57_wb_clk_i _02323_ _00619_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13848_ net1179 net1067 net3181 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[9\]
+ sky130_fd_sc_hd__and3b_1
X_17957__1472 vssd1 vssd1 vccd1 vccd1 _17957__1472/HI net1472 sky130_fd_sc_hd__conb_1
XFILLER_0_130_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12476__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16567_ clknet_leaf_158_wb_clk_i net830 _00550_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.ihit
+ sky130_fd_sc_hd__dfrtp_2
X_13779_ net1184 _04163_ vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__nand2_1
XANTENNA__14257__A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15518_ net1350 vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__inv_2
X_16498_ clknet_leaf_141_wb_clk_i _02252_ _00481_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15449_ net1237 vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10007__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1056 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09412__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_3_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold403 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[2\] vssd1 vssd1 vccd1 vccd1 net1938
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17119_ clknet_leaf_42_wb_clk_i _02806_ _01102_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold414 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[5\] vssd1 vssd1 vccd1 vccd1 net1949
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold425 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1960 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08620__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold436 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1971 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold447 _02151_ vssd1 vssd1 vccd1 vccd1 net1982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[13\] vssd1 vssd1 vccd1 vccd1
+ net1993 sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2004 sky130_fd_sc_hd__dlygate4sd3_1
X_09941_ _06280_ vssd1 vssd1 vccd1 vccd1 _06281_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_74_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout905 net906 vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__buf_2
XANTENNA__08421__C net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout916 _04779_ vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__buf_4
Xfanout927 net928 vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_146_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[12\] net798 net758 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06212_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_146_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout938 _04762_ vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__buf_4
Xfanout949 net950 vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ net1105 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[1\] net931 vssd1
+ vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__and3_1
Xhold1103 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1114 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2649 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout287_A _07896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_7__f_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_7__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1125 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2660 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1136 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2671 sky130_fd_sc_hd__dlygate4sd3_1
X_08754_ net1012 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[4\] net905 vssd1
+ vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__and3_1
Xhold1147 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[99\] vssd1 vssd1 vccd1 vccd1
+ net2682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1158 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2693 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09479__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1169 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2704 sky130_fd_sc_hd__dlygate4sd3_1
X_08685_ net1086 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[7\] net914 vssd1
+ vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout454_A _07957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12894__B net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12386__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09306_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[22\] net654 _05628_
+ _05642_ _05643_ vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_36_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10797__A1 _05963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09651__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09237_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[21\] net692 net660 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__a22o_1
XANTENNA__11303__B _05116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1151_X net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout507_X net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09939__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09168_ net1017 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[16\] net889 vssd1
+ vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__and3_1
XANTENNA__10549__A1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout990_A net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08119_ _04483_ team_01_WB.instance_to_wrap.cpu.f0.num\[10\] team_01_WB.instance_to_wrap.cpu.f0.num\[5\]
+ _04488_ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_107_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09099_ net1011 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[13\] net897 vssd1
+ vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__and3_1
XANTENNA__08611__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11130_ _06920_ _07216_ _07228_ _06928_ _07070_ vssd1 vssd1 vccd1 vccd1 _07470_ sky130_fd_sc_hd__a221o_1
Xhold970 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2505 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout876_X net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold981 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2516 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11061_ _05042_ _06438_ _07381_ _07399_ vssd1 vssd1 vccd1 vccd1 _07401_ sky130_fd_sc_hd__a2bb2o_1
Xhold992 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2527 sky130_fd_sc_hd__dlygate4sd3_1
X_10012_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[1\] _04634_ net795 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06352_ sky130_fd_sc_hd__a22o_1
X_14820_ net1220 vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__inv_2
XANTENNA__10222__X _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10589__B _06928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input15_A DAT_I[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11277__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14751_ net1189 vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__inv_2
XANTENNA__09162__C net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11963_ net3102 net216 net473 vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__mux2_1
XANTENNA__13671__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13702_ team_01_WB.instance_to_wrap.cpu.c0.count\[7\] _04103_ vssd1 vssd1 vccd1 vccd1
+ _04122_ sky130_fd_sc_hd__or2_1
X_17470_ clknet_leaf_80_wb_clk_i _03157_ _01453_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10914_ net341 net340 _06526_ net339 net550 net539 vssd1 vssd1 vccd1 vccd1 _07254_
+ sky130_fd_sc_hd__mux4_1
X_14682_ net1224 vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__inv_2
X_11894_ net2214 net221 net479 vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16421_ clknet_leaf_139_wb_clk_i _02175_ _00404_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10845_ _06921_ _06965_ vssd1 vssd1 vccd1 vccd1 _07185_ sky130_fd_sc_hd__or2_2
X_13633_ net186 _04069_ _04070_ net725 vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12296__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10237__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11434__C1 _07699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16352_ clknet_leaf_98_wb_clk_i _02106_ _00335_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[75\]
+ sky130_fd_sc_hd__dfrtp_1
X_10776_ _06641_ _06675_ _07114_ vssd1 vssd1 vccd1 vccd1 _07116_ sky130_fd_sc_hd__nand3_1
X_13564_ net185 _04011_ _04012_ net723 vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__a211o_1
XANTENNA__08075__A team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10788__A1 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09642__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15303_ net1389 vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16065__Q team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12515_ net3077 net298 net410 vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__mux2_1
XANTENNA__10892__X _07232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13495_ net196 net192 _07822_ net642 vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__o211a_1
XANTENNA__08850__B1 _05188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16283_ clknet_leaf_125_wb_clk_i _02037_ _00266_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13726__A1 net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12446_ net3096 net280 net418 vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15234_ net1320 vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08803__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12377_ net3045 net286 net425 vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__mux2_1
X_15165_ net1313 vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11328_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[4\] _07659_ vssd1 vssd1 vccd1
+ vccd1 _07662_ sky130_fd_sc_hd__nand2b_1
X_14116_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[62\] _04258_ _04263_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[126\]
+ _04401_ vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__a221o_1
X_15096_ net1215 vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11259_ _06935_ _07281_ _07597_ _07598_ vssd1 vssd1 vccd1 vccd1 _07599_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_52_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14047_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[11\] _04226_ _04244_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[99\]
+ _04335_ vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__a221o_1
XANTENNA__18012__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09634__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17806_ clknet_leaf_99_wb_clk_i _03482_ _01746_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[76\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15998_ net1408 vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_141_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17737_ clknet_leaf_116_wb_clk_i _03413_ _01677_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14949_ net1286 vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__inv_2
XANTENNA__10476__B1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08470_ net1119 net1125 net1122 net1116 vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__and4bb_4
X_17668_ clknet_leaf_158_wb_clk_i _03353_ _01609_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16619_ clknet_leaf_10_wb_clk_i _02306_ _00602_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_17599_ clknet_leaf_86_wb_clk_i _03286_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10719__S net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12768__A2 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09022_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[9\] net893 vssd1
+ vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__and3_1
XFILLER_0_143_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08713__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold200 net87 vssd1 vssd1 vccd1 vccd1 net1735 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13193__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold211 team_01_WB.instance_to_wrap.a1.ADR_I\[1\] vssd1 vssd1 vccd1 vccd1 net1746
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout202_A _07858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08432__B net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold222 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[120\] vssd1 vssd1 vccd1 vccd1
+ net1757 sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 team_01_WB.instance_to_wrap.cpu.f0.write_data\[3\] vssd1 vssd1 vccd1 vccd1
+ net1768 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1779 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold255 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1790 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12940__A2 _07757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold266 _02152_ vssd1 vssd1 vccd1 vccd1 net1801 sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1812 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[6\] vssd1 vssd1 vccd1 vccd1
+ net1823 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout702 _04758_ vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__buf_4
X_09924_ net1153 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[4\] net949 vssd1
+ vssd1 vccd1 vccd1 _06264_ sky130_fd_sc_hd__and3_1
Xhold299 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[19\] vssd1 vssd1 vccd1 vccd1 net1834
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout713 net714 vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12522__X _03565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1111_A net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout724 net728 vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1209_A net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout735 net736 vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__clkbuf_8
Xfanout746 net748 vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__clkbuf_8
X_09855_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[12\] net780 net753 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06195_ sky130_fd_sc_hd__a22o_1
Xfanout757 _04675_ vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__clkbuf_8
XANTENNA_input7_A DAT_I[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout768 _04672_ vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__buf_6
XANTENNA__10703__A1 _07042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout779 net781 vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__buf_6
XFILLER_0_147_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout669_A net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08806_ net1010 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[0\] net888 vssd1
+ vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__and3_1
X_09786_ net770 _06119_ _06122_ _06125_ vssd1 vssd1 vccd1 vccd1 _06126_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_134_Right_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08737_ net1017 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[4\] net922 vssd1
+ vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout836_A _03737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout457_X net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15281__A net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08668_ net1006 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[7\] net891 vssd1
+ vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__and3_1
XANTENNA__08447__X _04787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09872__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout624_X net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08599_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[15\] net669 _04937_ _04938_
+ vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__a211o_1
XFILLER_0_113_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10219__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16878__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10630_ net533 net503 vssd1 vssd1 vccd1 vccd1 _06970_ sky130_fd_sc_hd__nand2_1
XANTENNA__12759__A2 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10561_ _04736_ _04738_ vssd1 vssd1 vccd1 vccd1 _06901_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12844__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12300_ net2057 net203 net431 vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13280_ _03754_ _03768_ _04621_ vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10492_ net1131 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[31\] net956
+ vssd1 vssd1 vccd1 vccd1 _06832_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout993_X net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12231_ net2631 net248 net441 vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__mux2_1
XANTENNA__13184__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08342__B net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12931__A2 _07757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12162_ net2505 net210 net447 vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09157__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17956__1471 vssd1 vssd1 vccd1 vccd1 _17956__1471/HI net1471 sky130_fd_sc_hd__conb_1
XFILLER_0_20_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10942__A1 _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11113_ _06947_ _06951_ vssd1 vssd1 vccd1 vccd1 _07453_ sky130_fd_sc_hd__nor2_1
X_16970_ clknet_leaf_11_wb_clk_i _02657_ _00953_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_12093_ net2495 net223 net455 vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__mux2_1
X_11044_ _07382_ _07383_ vssd1 vssd1 vccd1 vccd1 _07384_ sky130_fd_sc_hd__nand2b_1
X_15921_ net1402 vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__inv_2
XANTENNA__11498__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08363__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15852_ net1334 vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__inv_2
XANTENNA__10170__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14803_ net1392 vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__inv_2
X_15783_ net1203 vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12995_ net2910 net2682 net861 vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__mux2_1
XANTENNA__11923__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17522_ clknet_leaf_113_wb_clk_i _03209_ _01505_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_14734_ net1211 vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__inv_2
X_11946_ net2886 net227 net475 vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09863__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17453_ clknet_leaf_67_wb_clk_i _03140_ _01436_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_14665_ net1228 vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__inv_2
X_11877_ net1885 net260 net485 vssd1 vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16404_ clknet_leaf_97_wb_clk_i net1889 _00387_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[127\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09076__A0 _05380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13616_ net186 _04055_ _04056_ net726 vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__a211o_1
X_17384_ clknet_leaf_62_wb_clk_i _03071_ _01367_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10828_ _07060_ _07100_ net327 _07082_ vssd1 vssd1 vccd1 vccd1 _07168_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_45_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14596_ net1362 vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__inv_2
XANTENNA__09615__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16335_ clknet_leaf_91_wb_clk_i net2223 _00318_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13547_ net185 _03997_ _03998_ net723 vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__a211o_1
XFILLER_0_137_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10759_ net532 _06935_ vssd1 vssd1 vccd1 vccd1 _07099_ sky130_fd_sc_hd__nor2_2
XANTENNA__18007__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09188__X _05528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09629__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16266_ clknet_leaf_151_wb_clk_i net1574 _00254_ vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13478_ _03934_ _03936_ _03938_ vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__or3_1
XANTENNA__17619__Q team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_18005_ net635 vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15217_ net1425 vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__inv_2
X_12429_ net1988 net246 net417 vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_93_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16197_ clknet_leaf_1_wb_clk_i _01957_ _00185_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_93_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10918__D1 _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13580__C1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15148_ net1259 vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10933__A1 _06912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15366__A net1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07970_ net1068 vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__inv_2
X_15079_ net1395 vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__inv_2
XANTENNA__08354__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09640_ net1135 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[23\] net972
+ vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_109_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_109_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09571_ net1149 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[25\] net977
+ vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_69_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11833__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08522_ net1078 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[18\] net883
+ vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__and3_1
XFILLER_0_132_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08453_ net1117 net1124 net1126 net1120 vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__and4bb_4
XFILLER_0_93_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08384_ net726 net719 vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14060__B1 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08814__B1 net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12664__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1061_A team_01_WB.instance_to_wrap.cpu.RU0.state\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout417_A _03562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire961_X net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10621__B1 _06960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1159_A net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09539__A net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09005_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[9\] net912 vssd1
+ vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13166__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10924__A1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout786_A _04659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09790__A1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08593__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14180__A net1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout510 _05996_ vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1114_X net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout521 _05260_ vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__buf_2
X_09907_ _06234_ _06235_ _06245_ _06246_ vssd1 vssd1 vccd1 vccd1 _06247_ sky130_fd_sc_hd__or4_1
Xfanout532 _05222_ vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__clkbuf_2
Xfanout543 net545 vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__clkbuf_4
Xfanout554 _05115_ vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__buf_2
XANTENNA_fanout953_A _04662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09705__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout565 net566 vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__buf_2
Xfanout576 _07792_ vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__buf_1
X_09838_ _06167_ _06170_ _06172_ _06177_ vssd1 vssd1 vccd1 vccd1 _06178_ sky130_fd_sc_hd__or4_1
Xfanout587 _04517_ vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__buf_2
Xfanout598 net599 vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__buf_4
XANTENNA__10152__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout741_X net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12839__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09769_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[15\] net802 net753 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout839_X net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11800_ net2078 net205 net491 vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__mux2_1
X_12780_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[16\] _07541_ net1034 vssd1 vssd1
+ vccd1 vccd1 _03615_ sky130_fd_sc_hd__mux2_1
X_11731_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[5\] net716 vssd1 vssd1 vccd1
+ vccd1 _07922_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14450_ net1204 vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_25_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[19\] _07135_ net713 vssd1 vssd1
+ vccd1 vccd1 _07867_ sky130_fd_sc_hd__mux2_1
XANTENNA__14051__B1 _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13401_ _03860_ _03861_ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_64_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10613_ _06951_ _06952_ vssd1 vssd1 vccd1 vccd1 _06953_ sky130_fd_sc_hd__nor2_1
XANTENNA__12574__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10883__A _05566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11593_ _07809_ vssd1 vssd1 vccd1 vccd1 _07810_ sky130_fd_sc_hd__inv_2
X_14381_ net1193 vssd1 vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16120_ clknet_leaf_135_wb_clk_i _01895_ _00108_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[27\]
+ sky130_fd_sc_hd__dfrtp_4
X_13332_ net564 _07702_ _03808_ net587 vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__a22o_1
X_10544_ _05805_ _05807_ _05835_ net561 vssd1 vssd1 vccd1 vccd1 _06884_ sky130_fd_sc_hd__a31o_1
Xwire966 net967 vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13157__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16051_ clknet_leaf_150_wb_clk_i _01844_ _00039_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_13263_ net1068 _03754_ team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1 vccd1
+ vccd1 _03755_ sky130_fd_sc_hd__o21ai_1
X_10475_ net504 _06780_ vssd1 vssd1 vccd1 vccd1 _06815_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_31_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15002_ net1371 vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__inv_2
X_12214_ net1879 net300 net444 vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12904__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13194_ net15 net837 net630 net3006 vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__a22o_1
XANTENNA__08033__B2 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10915__A1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11918__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_7_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12145_ net2885 net227 net451 vssd1 vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__mux2_1
XANTENNA__10391__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13314__C1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09184__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12076_ net1836 net258 net462 vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__mux2_1
X_16953_ clknet_leaf_102_wb_clk_i _02640_ _00936_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11027_ _05491_ _06158_ vssd1 vssd1 vccd1 vccd1 _07367_ sky130_fd_sc_hd__xor2_1
X_15904_ net1399 vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__inv_2
X_16884_ clknet_leaf_66_wb_clk_i _02571_ _00867_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10143__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15835_ net1331 vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__inv_2
XANTENNA__11576__A_N team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15766_ net1199 vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__inv_2
XANTENNA__13093__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08528__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12978_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[108\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[116\]
+ net860 vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__mux2_1
XANTENNA__09836__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17505_ clknet_leaf_54_wb_clk_i _03192_ _01488_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_38_wb_clk_i_X clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14717_ net1186 vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11929_ net2770 net214 net475 vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__mux2_1
X_15697_ net1395 vssd1 vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10496__C net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17436_ clknet_leaf_57_wb_clk_i _03123_ _01419_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_14648_ net1253 vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_70_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14042__B1 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_17 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_28 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12484__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17367_ clknet_leaf_15_wb_clk_i _03054_ _01350_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_39 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14579_ net1427 vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_60_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16318_ clknet_leaf_93_wb_clk_i _02072_ _00301_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08272__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17298_ clknet_leaf_110_wb_clk_i _02985_ _01281_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16249_ clknet_leaf_152_wb_clk_i net1635 _00237_ vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11159__A1 _06928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11159__B2 _06920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__buf_2
XANTENNA__13553__C1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__buf_2
Xoutput124 net124 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput135 net135 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__buf_2
Xoutput146 net146 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
Xoutput157 net157 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
XANTENNA__11828__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput168 net168 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__clkbuf_4
Xoutput179 net636 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire921_A _04775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11331__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09623_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] net626 _05961_ _05962_
+ vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_108_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13608__B1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12659__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09554_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[28\] net815 net737 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__a22o_1
XANTENNA__09827__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08438__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08505_ _04717_ _04752_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1 vssd1
+ vccd1 vccd1 _04845_ sky130_fd_sc_hd__o21a_1
XANTENNA__12869__B1_N net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12831__A1 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09485_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[30\] net665 net656 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__a22o_1
XANTENNA__12831__B2 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout534_A _05190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17955__1470 vssd1 vssd1 vccd1 vccd1 _17955__1470/HI net1470 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_156_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08436_ net1024 net919 vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__and2_2
Xclkbuf_leaf_77_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__14033__B1 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13998__B team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08367_ _04706_ vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__inv_2
XANTENNA__12394__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout701_A _04758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08298_ net1164 net1167 net1158 net1161 vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__and4bb_1
XANTENNA__09460__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13139__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10260_ _06133_ _06162_ _06165_ _06599_ _06132_ vssd1 vssd1 vccd1 vccd1 _06600_ sky130_fd_sc_hd__o221a_1
XFILLER_0_42_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08460__X _04800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout691_X net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout789_X net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ _06528_ _06529_ _06526_ vssd1 vssd1 vccd1 vccd1 _06531_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_115_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1305 net1306 vssd1 vssd1 vccd1 vccd1 net1305 sky130_fd_sc_hd__buf_4
Xfanout1316 net1321 vssd1 vssd1 vccd1 vccd1 net1316 sky130_fd_sc_hd__buf_4
Xfanout1327 net1332 vssd1 vssd1 vccd1 vccd1 net1327 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout340 _06495_ vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__clkbuf_4
Xfanout1338 net1344 vssd1 vssd1 vccd1 vccd1 net1338 sky130_fd_sc_hd__buf_4
XANTENNA_fanout956_X net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout351 _03742_ vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1349 net1369 vssd1 vssd1 vccd1 vccd1 net1349 sky130_fd_sc_hd__buf_2
XANTENNA__15734__A net1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout362 _03580_ vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__clkbuf_4
X_13950_ _04223_ _04227_ vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__nand2_2
Xfanout373 _06188_ vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__clkbuf_4
Xfanout384 _03570_ vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__buf_4
Xfanout395 _03567_ vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__clkbuf_8
X_12901_ net360 _03675_ net1036 vssd1 vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09732__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13881_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[3\] _04187_ vssd1 vssd1 vccd1
+ vccd1 _04188_ sky130_fd_sc_hd__and2_1
XANTENNA__12569__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13254__A team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15620_ net1222 vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__inv_2
X_12832_ net1620 net639 net606 _03650_ vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15551_ net1311 vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__inv_2
X_12763_ net1691 net638 net606 _03603_ vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14502_ net1354 vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__inv_2
X_11714_ net1963 net281 net500 vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15482_ net1372 vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__inv_2
XANTENNA__14024__B1 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12694_ net2503 net206 net385 vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17221_ clknet_leaf_53_wb_clk_i _02908_ _01204_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14433_ net1306 vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__inv_2
X_11645_ _07817_ _07853_ vssd1 vssd1 vccd1 vccd1 _07854_ sky130_fd_sc_hd__and2b_1
XFILLER_0_86_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12157__X _07958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17152_ clknet_leaf_47_wb_clk_i _02839_ _01135_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09179__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput15 DAT_I[21] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
X_14364_ net1206 vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_154_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xinput26 DAT_I[31] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
X_11576_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\]
+ vssd1 vssd1 vccd1 vccd1 _07793_ sky130_fd_sc_hd__and2b_1
Xinput37 gpio_in[19] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_1
XFILLER_0_24_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16073__Q team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16103_ clknet_leaf_127_wb_clk_i _01878_ _00091_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[10\]
+ sky130_fd_sc_hd__dfrtp_2
Xinput48 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_1
X_13315_ _04475_ _07706_ vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__nand2_1
Xinput59 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08514__C net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17083_ clknet_leaf_74_wb_clk_i _02770_ _01066_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10527_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[31\] net696 net672 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[31\]
+ _06866_ vssd1 vssd1 vccd1 vccd1 _06867_ sky130_fd_sc_hd__a221o_1
X_14295_ net1328 vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__inv_2
X_16034_ clknet_leaf_135_wb_clk_i _01828_ _00028_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13246_ net2702 net354 net350 team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1
+ vccd1 vccd1 _01904_ sky130_fd_sc_hd__a22o_1
X_10458_ _06795_ _06796_ _06797_ vssd1 vssd1 vccd1 vccd1 _06798_ sky130_fd_sc_hd__or3_1
XFILLER_0_149_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12889__A1 _05704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11648__S net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13429__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10389_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[16\] net816 _06727_
+ _06728_ vssd1 vssd1 vccd1 vccd1 _06729_ sky130_fd_sc_hd__a211o_1
X_13177_ net1 _03732_ vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__nand2_1
X_12128_ net2228 net215 net451 vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__mux2_1
X_17985_ net1500 vssd1 vssd1 vccd1 vccd1 la_data_out[27] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_36_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09345__C net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16936_ clknet_leaf_62_wb_clk_i _02623_ _00919_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_12059_ net2153 net188 net459 vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__mux2_1
XANTENNA__10116__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11313__A1 _04504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12479__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16867_ clknet_leaf_27_wb_clk_i _02554_ _00850_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_15818_ net1190 vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__inv_2
X_16798_ clknet_leaf_84_wb_clk_i _02485_ _00781_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09080__C net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15749_ net1341 vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_103_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12813__B2 _03637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09270_ _05604_ _05605_ _05607_ _05609_ vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_62_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14015__B1 _04265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08221_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[60\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[52\]
+ net1050 vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17419_ clknet_leaf_7_wb_clk_i _03106_ _01402_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09089__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08152_ net829 net566 vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_151_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09442__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08424__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08083_ net1818 net569 _04525_ _04556_ vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_124_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_124_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10355__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1024_A net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08440__B net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08985_ net1007 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[8\] net929 vssd1
+ vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout484_A _07948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10107__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout651_A _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12389__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout749_A _04680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09606_ net1146 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[24\] net952
+ vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__and3_1
XANTENNA__08720__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11068__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09537_ net996 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[28\] net979 vssd1
+ vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__and3_1
XFILLER_0_149_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12804__A1 _07290_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1181_X net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout916_A _04779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14006__B1 _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09468_ net561 _05805_ _05807_ vssd1 vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__o21a_1
XFILLER_0_109_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09681__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08419_ net1116 net1125 net1122 net1119 vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__and4bb_4
XANTENNA_fanout704_X net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09399_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[27\] net690 net665 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11430_ team_01_WB.instance_to_wrap.cpu.f0.i\[11\] _07676_ net610 team_01_WB.instance_to_wrap.cpu.f0.i\[12\]
+ vssd1 vssd1 vccd1 vccd1 _07740_ sky130_fd_sc_hd__a31o_1
XFILLER_0_151_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09433__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11361_ team_01_WB.instance_to_wrap.cpu.f0.i\[16\] team_01_WB.instance_to_wrap.cpu.f0.i\[15\]
+ _07689_ vssd1 vssd1 vccd1 vccd1 _07690_ sky130_fd_sc_hd__and3_1
XANTENNA__11240__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14055__D _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12852__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_886 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14633__A net1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13517__C1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13100_ net52 net51 net54 net53 vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__or4_1
X_10312_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[18\] net782 net739 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06652_ sky130_fd_sc_hd__a22o_1
X_11292_ _07628_ net1169 _07631_ vssd1 vssd1 vccd1 vccd1 _07632_ sky130_fd_sc_hd__mux2_1
X_14080_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[100\] _04244_ _04255_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[116\]
+ vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__a22o_1
XANTENNA__08631__A team_01_WB.instance_to_wrap.cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_120_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08539__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10243_ _06576_ _06577_ _06578_ _06582_ vssd1 vssd1 vccd1 vccd1 _06583_ sky130_fd_sc_hd__or4_1
X_13031_ net2757 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[63\] net856 vssd1 vssd1
+ vccd1 vccd1 _02094_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10174_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[10\] net813 net758 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06514_ sky130_fd_sc_hd__a22o_1
Xfanout1102 net1103 vssd1 vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input45_A wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1113 net1114 vssd1 vssd1 vccd1 vccd1 net1113 sky130_fd_sc_hd__clkbuf_2
Xfanout1124 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[21\] vssd1 vssd1 vccd1 vccd1
+ net1124 sky130_fd_sc_hd__buf_2
Xfanout1135 net1141 vssd1 vssd1 vccd1 vccd1 net1135 sky130_fd_sc_hd__buf_2
X_17770_ clknet_leaf_123_wb_clk_i _03446_ _01710_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[40\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1146 net1151 vssd1 vssd1 vccd1 vccd1 net1146 sky130_fd_sc_hd__buf_1
X_14982_ net1405 vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__inv_2
XANTENNA__13296__A1 _07650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1157 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[19\] vssd1 vssd1 vccd1 vccd1
+ net1157 sky130_fd_sc_hd__buf_2
Xfanout1168 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[15\] vssd1 vssd1 vccd1 vccd1
+ net1168 sky130_fd_sc_hd__buf_2
XANTENNA__10104__C net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1179 net1180 vssd1 vssd1 vccd1 vccd1 net1179 sky130_fd_sc_hd__clkbuf_2
Xfanout192 _07634_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__clkbuf_4
X_16721_ clknet_leaf_116_wb_clk_i _02408_ _00704_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13933_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__nand2_8
XANTENNA__12299__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16652_ clknet_leaf_16_wb_clk_i _02339_ _00635_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13864_ net1178 net1064 net1643 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[25\]
+ sky130_fd_sc_hd__and3b_1
XANTENNA__10401__A net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15603_ net1383 vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_83_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16068__Q team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12815_ net1038 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[5\] vssd1 vssd1 vccd1
+ vccd1 _03639_ sky130_fd_sc_hd__or2_1
XANTENNA__08509__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16583_ clknet_leaf_106_wb_clk_i _02270_ _00566_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13795_ _04165_ _04176_ vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11931__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15534_ net1291 vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__inv_2
X_12746_ net1745 net639 net607 _03591_ vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08806__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15465_ net1293 vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__inv_2
XANTENNA__08119__A1_N _04483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11325__B1_N team_01_WB.instance_to_wrap.cpu.DM0.data_i\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12677_ net2280 net282 net390 vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__mux2_1
X_17204_ clknet_leaf_23_wb_clk_i _02891_ _01187_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_14416_ net1308 vssd1 vssd1 vccd1 vccd1 _00210_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11628_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] _07818_ vssd1 vssd1
+ vccd1 vccd1 _07840_ sky130_fd_sc_hd__nor2_1
X_15396_ net1220 vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__inv_2
XANTENNA__09424__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09975__A1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17135_ clknet_leaf_31_wb_clk_i _02822_ _01118_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13771__A2 _04152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14347_ net1333 vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__inv_2
XANTENNA__09975__B2 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap304 _07188_ vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__clkbuf_2
X_11559_ _07787_ _07788_ vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__nor2_1
XANTENNA__18015__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire582 _06096_ vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10585__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold607 net113 vssd1 vssd1 vccd1 vccd1 net2142 sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2153 sky130_fd_sc_hd__dlygate4sd3_1
Xhold629 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2164 sky130_fd_sc_hd__dlygate4sd3_1
X_17066_ clknet_leaf_32_wb_clk_i _02753_ _01049_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_14278_ net1340 vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_38_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17627__Q team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09727__A1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16017_ net1329 vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__inv_2
X_13229_ net2752 net352 net348 team_01_WB.instance_to_wrap.cpu.f0.i\[21\] vssd1 vssd1
+ vccd1 vccd1 _01921_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12731__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11534__B2 net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08950__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1307 _02133_ vssd1 vssd1 vccd1 vccd1 net2842 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_4_6__f_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_6__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xhold1318 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2853 sky130_fd_sc_hd__dlygate4sd3_1
X_08770_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[4\] net704 _05104_ _05109_
+ vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__o22a_4
X_17968_ net1483 vssd1 vssd1 vccd1 vccd1 la_data_out[10] sky130_fd_sc_hd__buf_2
XFILLER_0_97_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1329 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[73\] vssd1 vssd1 vccd1 vccd1
+ net2864 sky130_fd_sc_hd__dlygate4sd3_1
X_16919_ clknet_leaf_16_wb_clk_i _02606_ _00902_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_144_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17899_ net1434 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_105_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08702__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12002__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12798__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11841__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09322_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[24\] net681 net669 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08716__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09253_ net600 _05592_ vssd1 vssd1 vccd1 vccd1 _05593_ sky130_fd_sc_hd__or2_2
XANTENNA__11470__B1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout232_A _07884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08204_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[77\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[69\]
+ net1050 vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__mux2_1
X_09184_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[16\] net879
+ vssd1 vssd1 vccd1 vccd1 _05524_ sky130_fd_sc_hd__and3_1
XFILLER_0_146_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08135_ _04489_ team_01_WB.instance_to_wrap.cpu.f0.num\[0\] team_01_WB.instance_to_wrap.cpu.f0.num\[19\]
+ _04475_ vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_16_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12672__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1141_A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10576__A2 _06882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08066_ _04512_ _04529_ _04539_ vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout699_A _04760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13514__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1406_A net1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11525__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout866_A net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout487_X net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08968_ net1007 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[8\] net900 vssd1
+ vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_125_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08899_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[2\] net889 vssd1
+ vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout654_X net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_3_Left_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10930_ _06469_ _06472_ _06568_ vssd1 vssd1 vccd1 vccd1 _07270_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_92_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_98_558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout821_X net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10861_ net522 _07123_ _07149_ _06957_ vssd1 vssd1 vccd1 vccd1 _07201_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_21_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12847__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14628__A net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout919_X net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12789__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12600_ net2673 net271 net395 vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13580_ net198 net194 _07879_ net644 vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10792_ net515 _06897_ _07120_ vssd1 vssd1 vccd1 vccd1 _07132_ sky130_fd_sc_hd__o21a_1
XANTENNA__13450__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12531_ net2061 net205 net403 vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08345__B net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11052__A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15250_ net1292 vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__inv_2
XANTENNA__09406__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12462_ net2806 net246 net413 vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__mux2_1
X_18013__1511 vssd1 vssd1 vccd1 vccd1 _18013__1511/HI net1511 sky130_fd_sc_hd__conb_1
XFILLER_0_53_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14201_ net1695 vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__clkbuf_1
X_11413_ _07693_ _07729_ vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__nor2_1
X_15181_ net1268 vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__inv_2
XANTENNA__12582__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14363__A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11202__D _07541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12393_ net2837 net220 net421 vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14132_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[71\] _04247_ _04249_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__a22o_1
X_11344_ team_01_WB.instance_to_wrap.cpu.f0.i\[2\] team_01_WB.instance_to_wrap.cpu.f0.i\[1\]
+ _07671_ vssd1 vssd1 vccd1 vccd1 _07673_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14063_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[99\] _04254_ _04263_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[123\]
+ vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__a22o_1
X_11275_ _07038_ _07100_ net327 _07029_ vssd1 vssd1 vccd1 vccd1 _07615_ sky130_fd_sc_hd__a22o_1
XANTENNA__11516__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10319__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_148_Right_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13014_ net2801 net2794 net857 vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__mux2_1
X_10226_ _06562_ _06565_ vssd1 vssd1 vccd1 vccd1 _06566_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_33_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11926__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10157_ net560 _04970_ _05378_ vssd1 vssd1 vccd1 vccd1 _06497_ sky130_fd_sc_hd__or3_1
X_17822_ clknet_leaf_119_wb_clk_i _03498_ _01762_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[92\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__13269__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 team_01_WB.instance_to_wrap.cpu.RU0.state\[1\] vssd1 vssd1 vccd1 vccd1 net1539
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09192__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10088_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[7\] net760 _06417_ _06420_
+ net769 vssd1 vssd1 vccd1 vccd1 _06428_ sky130_fd_sc_hd__a2111o_1
X_14965_ net1282 vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_50_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17753_ clknet_leaf_121_wb_clk_i net2592 _01693_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16704_ clknet_leaf_48_wb_clk_i _02391_ _00687_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13916_ _04142_ _04207_ vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__and2_1
X_17684_ clknet_leaf_129_wb_clk_i _03368_ _01625_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10131__A net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14896_ net1270 vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_18_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16635_ clknet_leaf_69_wb_clk_i _02322_ _00618_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13847_ net1181 team_01_WB.instance_to_wrap.cpu.RU0.state\[4\] team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[8\]
+ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[8\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_58_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11661__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13442__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16566_ clknet_leaf_157_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_dhit _00549_
+ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.dhit sky130_fd_sc_hd__dfrtp_4
XFILLER_0_128_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13778_ team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[2\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[2\]
+ net605 vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__mux2_1
XANTENNA__09645__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_0_0_wb_clk_i_X clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15517_ net1313 vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__inv_2
X_12729_ _03575_ _03578_ vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16497_ clknet_leaf_151_wb_clk_i _02251_ _00480_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13992__A2 _04245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15448_ net1212 vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13744__A2 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12492__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15379_ net1383 vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17118_ clknet_leaf_82_wb_clk_i _02805_ _01101_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold404 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1939 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold415 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold426 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1961 sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1972 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold448 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[17\] vssd1 vssd1 vccd1 vccd1
+ net1983 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14154__C1 net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold459 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1994 sky130_fd_sc_hd__dlygate4sd3_1
X_09940_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] net626 _06278_ _06279_
+ vssd1 vssd1 vccd1 vccd1 _06280_ sky130_fd_sc_hd__a22o_4
X_17049_ clknet_leaf_103_wb_clk_i _02736_ _01032_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09654__X _05994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout906 _04785_ vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__clkbuf_8
X_09871_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[12\] net743 net735 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06211_ sky130_fd_sc_hd__a22o_1
Xfanout917 net918 vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_146_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout928 _04767_ vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__buf_4
Xfanout939 net940 vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_146_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11836__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08822_ net1022 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[1\] net942 vssd1
+ vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__and3_1
XANTENNA__10740__S net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10191__B1 _06526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1104 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2639 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1115 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2650 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1126 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[59\] vssd1 vssd1 vccd1 vccd1
+ net2661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2672 sky130_fd_sc_hd__dlygate4sd3_1
X_08753_ net1094 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[4\] net905 vssd1
+ vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__and3_1
XFILLER_0_139_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1148 team_01_WB.instance_to_wrap.cpu.f0.num\[14\] vssd1 vssd1 vccd1 vccd1 net2683
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09533__C net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1159 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[51\] vssd1 vssd1 vccd1 vccd1
+ net2694 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10041__A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08684_ net1086 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[7\] net888 vssd1
+ vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_120_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11691__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12667__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1091_A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout447_A _07958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08446__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09305_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[22\] net679 _05630_
+ _05636_ _05637_ vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11443__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_48_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13983__A2 _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10797__A2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09236_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[21\] net668 _05574_ _05575_
+ vssd1 vssd1 vccd1 vccd1 _05576_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_118_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13196__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09939__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13735__A2 _04574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout402_X net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09167_ net1091 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[16\] net882
+ vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09403__A3 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1144_X net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11600__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09277__A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08118_ net1069 _04495_ team_01_WB.instance_to_wrap.cpu.f0.num\[18\] _04476_ vssd1
+ vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__a22o_1
XANTENNA__08611__A1 net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09098_ net1011 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[13\] net934 vssd1
+ vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09708__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08049_ _04521_ team_01_WB.instance_to_wrap.cpu.K0.code\[3\] team_01_WB.instance_to_wrap.cpu.K0.code\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__or3b_2
XFILLER_0_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold960 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold971 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2506 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1409_X net1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold982 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2517 sky130_fd_sc_hd__dlygate4sd3_1
X_11060_ net372 _07380_ _05301_ vssd1 vssd1 vccd1 vccd1 _07400_ sky130_fd_sc_hd__nor3b_1
Xhold993 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2528 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout771_X net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout869_X net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12171__A1 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10011_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[1\] net751 net770 vssd1
+ vssd1 vccd1 vccd1 _06351_ sky130_fd_sc_hd__a21o_1
XANTENNA__08914__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10182__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_Left_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09443__C net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13120__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11047__A net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14750_ net1187 vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__inv_2
X_11962_ net3042 net219 net473 vssd1 vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__mux2_1
XANTENNA__09875__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13701_ _04106_ _04119_ _04121_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[9\]
+ sky130_fd_sc_hd__and3b_1
XANTENNA__09740__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10913_ _06596_ _07252_ vssd1 vssd1 vccd1 vccd1 _07253_ sky130_fd_sc_hd__xor2_1
XANTENNA__12577__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14681_ net1227 vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__inv_2
X_11893_ net2942 net188 net479 vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__mux2_1
XANTENNA__13262__A team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16420_ clknet_leaf_130_wb_clk_i _02174_ _00403_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13632_ net197 net193 _07911_ net643 vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__o211a_1
X_10844_ net338 _07016_ net328 _07183_ _07179_ vssd1 vssd1 vccd1 vccd1 _07184_ sky130_fd_sc_hd__a221o_1
XANTENNA__13423__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13423__B2 net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16351_ clknet_leaf_90_wb_clk_i net2780 _00334_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13563_ net196 net192 _07869_ net642 vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__o211a_1
X_10775_ _06675_ _07114_ _06641_ vssd1 vssd1 vccd1 vccd1 _07115_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15302_ net1380 vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__inv_2
X_12514_ net1914 net276 net408 vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__mux2_1
X_16282_ clknet_leaf_116_wb_clk_i _02036_ _00265_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[5\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_57_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13494_ _03952_ _03954_ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08850__A1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13187__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15233_ net1279 vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__inv_2
X_12445_ net3017 net251 net418 vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15164_ net1243 vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__inv_2
X_12376_ net2136 net253 net424 vssd1 vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__mux2_1
X_14115_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[62\] _04260_ _04267_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__a22o_1
XANTENNA__08522__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11327_ _07661_ net2036 _07655_ vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__mux2_1
X_15095_ net1249 vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__inv_2
XANTENNA__09915__A _06250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14151__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14046_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[35\] _04221_ _04230_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[35\]
+ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__a22o_1
X_11258_ _06966_ _07278_ _06964_ vssd1 vssd1 vccd1 vccd1 _07598_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08366__B1 _04704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11656__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10209_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[8\] net819 net814 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _06549_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_66_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11189_ _06921_ _07527_ _07528_ _07185_ vssd1 vssd1 vccd1 vccd1 _07529_ sky130_fd_sc_hd__o211ai_1
X_17805_ clknet_leaf_95_wb_clk_i _03481_ _01745_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[75\]
+ sky130_fd_sc_hd__dfrtp_1
X_15997_ net1417 vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_141_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10499__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14948_ net1218 vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__inv_2
X_17736_ clknet_leaf_116_wb_clk_i _03412_ _01676_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09866__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10476__A1 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09330__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12487__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17667_ clknet_leaf_157_wb_clk_i _03352_ _01608_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17640__Q team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14879_ net1311 vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__inv_2
X_16618_ clknet_leaf_32_wb_clk_i _02305_ _00601_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_17598_ clknet_leaf_86_wb_clk_i _03285_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09618__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16549_ clknet_leaf_1_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[15\]
+ _00532_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_75_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09021_ net1095 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[9\] net925 vssd1
+ vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold201 _02018_ vssd1 vssd1 vccd1 vccd1 net1736 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold212 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1747 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold223 _03526_ vssd1 vssd1 vccd1 vccd1 net1758 sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1769 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold245 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1780 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold256 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[8\] vssd1 vssd1 vccd1 vccd1
+ net1791 sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 net82 vssd1 vssd1 vccd1 vccd1 net1802 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold278 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 net1813
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ net1153 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[4\] net971 vssd1
+ vssd1 vccd1 vccd1 _06263_ sky130_fd_sc_hd__and3_1
Xfanout703 _04758_ vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__buf_8
XANTENNA__14142__A2 _04236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold289 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1824 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout714 net717 vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_84_Left_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08357__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13853__A_N net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout725 net728 vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout397_A _03567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout736 _04687_ vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__buf_8
Xfanout747 net748 vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__clkbuf_4
X_09854_ _06192_ _06193_ vssd1 vssd1 vccd1 vccd1 _06194_ sky130_fd_sc_hd__nand2b_1
Xfanout758 _04675_ vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__clkbuf_4
Xfanout769 _04672_ vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1104_A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08805_ net1093 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[0\] net897 vssd1
+ vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__and3_1
X_09785_ _06109_ _06110_ _06123_ _06124_ vssd1 vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout564_A net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout185_X net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08736_ net602 _05074_ _05075_ vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__a21o_1
XANTENNA__13653__A1 _07639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10202__C net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09321__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08667_ net1006 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[7\] net914 vssd1
+ vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout731_A net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12397__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1094_X net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09609__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08598_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[15\] net686 net666 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_93_Left_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10560_ _04741_ _04743_ vssd1 vssd1 vccd1 vccd1 _06900_ sky130_fd_sc_hd__nand2_2
XFILLER_0_91_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08904__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09219_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[17\] net683 _05547_
+ _05548_ _05552_ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_20_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10491_ net1131 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[31\] net981
+ vssd1 vssd1 vccd1 vccd1 _06831_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_20_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12916__B1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12230_ net2225 net211 net439 vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout986_X net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08596__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12860__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12161_ net2783 net216 net449 vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10942__A2 _06707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11112_ net551 _06465_ _06946_ vssd1 vssd1 vccd1 vccd1 _07452_ sky130_fd_sc_hd__o21ba_1
XANTENNA__09735__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14133__A2 _04246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12092_ net1939 net189 net455 vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__mux2_1
Xhold790 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2325 sky130_fd_sc_hd__dlygate4sd3_1
X_11043_ _05076_ _06250_ vssd1 vssd1 vccd1 vccd1 _07383_ sky130_fd_sc_hd__nand2_1
X_15920_ net1401 vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__inv_2
X_15851_ net1334 vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__inv_2
XANTENNA__09173__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14802_ net1290 vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__inv_2
X_15782_ net1203 vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09848__B1 _06186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13644__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12994_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[92\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[100\]
+ net860 vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__mux2_1
XANTENNA__10887__Y _07227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1490 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net3025 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09470__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14733_ net1211 vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__inv_2
X_17521_ clknet_leaf_117_wb_clk_i _03208_ _01504_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09312__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11945_ net2379 net284 net478 vssd1 vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17452_ clknet_leaf_19_wb_clk_i _03139_ _01435_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_14664_ net1307 vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__inv_2
XANTENNA__12100__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11876_ net1997 net230 net485 vssd1 vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_60_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16403_ clknet_leaf_120_wb_clk_i net1876 _00386_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[126\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13615_ net199 net195 _07806_ _07899_ net644 vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__o2111a_1
XANTENNA__08517__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10827_ net369 _07165_ _07166_ net507 _05619_ vssd1 vssd1 vccd1 vccd1 _07167_ sky130_fd_sc_hd__o32a_1
XANTENNA__09076__A1 _05415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17383_ clknet_leaf_100_wb_clk_i _03070_ _01366_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_14595_ net1359 vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14816__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16334_ clknet_leaf_93_wb_clk_i net2445 _00317_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13546_ net196 net192 _07857_ net642 vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__o211a_1
X_10758_ _04844_ net331 _07094_ net369 _07097_ vssd1 vssd1 vccd1 vccd1 _07098_ sky130_fd_sc_hd__a221o_1
XFILLER_0_82_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16265_ clknet_leaf_151_wb_clk_i net1597 _00253_ vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__dfrtp_1
X_13477_ _04500_ _04842_ _03937_ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10689_ _07027_ _07028_ net519 vssd1 vssd1 vccd1 vccd1 _07029_ sky130_fd_sc_hd__mux2_1
X_18004_ net636 vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15216_ net1273 vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_134_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09379__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12428_ net2233 net210 net415 vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16196_ clknet_leaf_1_wb_clk_i _01956_ _00184_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_93_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14109__C1 net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15147_ net1424 vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__inv_2
XANTENNA__12770__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12359_ net2097 net221 net423 vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14124__A2 _04221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15078_ net1381 vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__inv_2
X_14029_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[2\] _04249_ _04259_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[18\]
+ _04318_ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__a221o_1
XANTENNA__09551__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09083__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09570_ net997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[25\] net955 vssd1
+ vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__and3_1
XANTENNA__09839__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13635__A1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08521_ net1081 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[18\] net935
+ vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__and3_1
X_17719_ clknet_leaf_156_wb_clk_i _00014_ _01660_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_69_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_149_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_149_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11415__A team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12010__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08452_ net1082 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[23\] net944
+ vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08383_ net1170 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[4\]
+ _04711_ vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__or4_1
XANTENNA__14726__A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08814__A1 _04708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10973__B net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10621__A1 _06886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout312_A _07931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08443__B net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09004_ net1013 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[9\] net917 vssd1
+ vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__and3_1
XANTENNA__11150__A _07476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12680__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10385__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08042__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1221_A net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_105_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10924__A2 _07263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1319_A net1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14115__A2 _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout681_A _04787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout500 net501 vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout779_A net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout511 _05963_ vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__clkbuf_4
X_09906_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[5\] net818 net751 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06246_ sky130_fd_sc_hd__a22o_1
Xfanout522 net527 vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11149__X _07489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout533 _05190_ vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10137__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout544 net545 vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__clkbuf_2
Xfanout555 net556 vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__buf_2
Xfanout566 _04620_ vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__clkbuf_2
X_09837_ _06173_ _06174_ _06175_ _06176_ vssd1 vssd1 vccd1 vccd1 _06177_ sky130_fd_sc_hd__or4_1
Xfanout577 net578 vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__buf_2
Xfanout588 net589 vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__buf_2
Xfanout599 _04755_ vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__clkbuf_4
XANTENNA__15292__A net1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09768_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[15\] net750 net740 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06108_ sky130_fd_sc_hd__a22o_1
XANTENNA__09290__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08719_ net1098 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[5\] net893 vssd1
+ vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__and3_1
X_09699_ net997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[21\] net955 vssd1
+ vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout734_X net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11730_ net1936 net296 net500 vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08337__C net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout901_X net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11661_ net2593 net271 net501 vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__mux2_1
XANTENNA__12855__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13400_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] net595 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10612_ net551 _06339_ vssd1 vssd1 vccd1 vccd1 _06952_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14380_ net1195 vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__inv_2
X_11592_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] _07808_ vssd1 vssd1
+ vccd1 vccd1 _07809_ sky130_fd_sc_hd__and2_1
XANTENNA__08634__A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10883__B _06707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_144_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_135_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13331_ _04479_ _07686_ _03743_ vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_148_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10543_ net503 _06882_ vssd1 vssd1 vccd1 vccd1 _06883_ sky130_fd_sc_hd__xor2_4
XANTENNA__11060__A net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16050_ clknet_leaf_148_wb_clk_i _01843_ _00038_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_13262_ team_01_WB.instance_to_wrap.cpu.f0.i\[26\] _03753_ vssd1 vssd1 vccd1 vccd1
+ _03754_ sky130_fd_sc_hd__or2_1
Xwire978 _04635_ vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__clkbuf_2
X_10474_ _06811_ _06813_ vssd1 vssd1 vccd1 vccd1 _06814_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09168__C net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15001_ net1238 vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__inv_2
X_12213_ net2401 net282 net446 vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__mux2_1
XANTENNA__12590__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13193_ net16 net835 net628 net1660 vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__o22a_1
XFILLER_0_32_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10915__A2 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12144_ net3118 net286 net453 vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__mux2_1
XANTENNA__14106__A2 _04230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09781__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16952_ clknet_leaf_49_wb_clk_i _02639_ _00935_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12075_ net2342 net231 net461 vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__mux2_1
XANTENNA__10679__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11026_ _04947_ net374 vssd1 vssd1 vccd1 vccd1 _07366_ sky130_fd_sc_hd__xor2_1
X_15903_ net1411 vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16883_ clknet_leaf_24_wb_clk_i _02570_ _00866_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11934__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15834_ net1331 vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__inv_2
XANTENNA__13617__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15765_ net1198 vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09631__C net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12977_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[109\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[117\]
+ net859 vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17504_ clknet_leaf_48_wb_clk_i _03191_ _01487_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_14716_ net1186 vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__inv_2
X_11928_ net2884 net218 net477 vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__mux2_1
X_15696_ net1271 vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17435_ clknet_leaf_70_wb_clk_i _03122_ _01418_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_14647_ net1314 vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__inv_2
X_11859_ net575 _07793_ _07946_ vssd1 vssd1 vccd1 vccd1 _07948_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_64_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14042__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_18 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_144_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_29 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14578_ net1366 vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__inv_2
X_17366_ clknet_leaf_30_wb_clk_i _03053_ _01349_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16534__Q team_01_WB.instance_to_wrap.cpu.DM0.data_i\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13529_ net187 _03982_ _03983_ net727 vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__a211o_1
X_16317_ clknet_leaf_120_wb_clk_i _02071_ _00300_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17297_ clknet_leaf_117_wb_clk_i _02984_ _01280_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_18003__1507 vssd1 vssd1 vccd1 vccd1 _18003__1507/HI net1507 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_132_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16248_ clknet_leaf_151_wb_clk_i net1631 _00236_ vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__buf_2
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__buf_2
X_16179_ clknet_leaf_7_wb_clk_i _01939_ _00167_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_110_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput125 net125 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__buf_2
XFILLER_0_140_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput136 net136 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__buf_2
XANTENNA__10906__A2 _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput147 net147 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_103_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput158 net158 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
XANTENNA__09772__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput169 net169 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12108__A1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08710__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12005__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10119__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10314__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09524__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11844__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09622_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[24\] net765 net624 vssd1
+ vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_108_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13608__A1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08719__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11619__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09553_ _05876_ _05890_ _05891_ _05892_ vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__or4_1
XFILLER_0_78_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09541__C _04640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout262_A _07880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08438__B net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08504_ net597 _04837_ _04843_ vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__o21a_2
XANTENNA__11145__A _05263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09484_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[30\] net646 _05812_
+ _05813_ _05815_ vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_148_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12831__A2 _07438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08435_ net1116 net1119 net1122 net1125 vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__nor4b_2
XTAP_TAPCELL_ROW_156_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12675__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1171_A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1269_A net1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08366_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] net625 _04704_ _04705_
+ vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__a22o_4
XANTENNA__08454__A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08297_ net991 net981 vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_46_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__17643__CLK clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout896_A net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10358__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10190_ _06526_ _06528_ _06529_ vssd1 vssd1 vccd1 vccd1 _06530_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout684_X net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1306 net1322 vssd1 vssd1 vccd1 vccd1 net1306 sky130_fd_sc_hd__buf_4
Xfanout1317 net1321 vssd1 vssd1 vccd1 vccd1 net1317 sky130_fd_sc_hd__buf_4
Xfanout330 _06924_ vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__clkbuf_4
Xfanout1328 net1332 vssd1 vssd1 vccd1 vccd1 net1328 sky130_fd_sc_hd__buf_4
Xfanout341 _06216_ vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__clkbuf_4
Xfanout1339 net1344 vssd1 vssd1 vccd1 vccd1 net1339 sky130_fd_sc_hd__clkbuf_4
Xfanout352 net353 vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__buf_2
XFILLER_0_100_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout363 _03580_ vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__buf_2
XANTENNA_fanout851_X net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout374 _06129_ vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__clkbuf_4
Xfanout385 _03570_ vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__buf_6
XANTENNA_fanout949_X net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout396 _03567_ vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__clkbuf_4
X_12900_ _05654_ net577 vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__nor2_1
XANTENNA__11754__S net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13880_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[2\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[1\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1 _04187_
+ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_21_Left_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12831_ net1033 _07438_ net362 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\]
+ net1060 vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__a32o_1
XFILLER_0_68_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08348__B net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15550_ net1321 vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__inv_2
X_12762_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] net1061 net362 _03602_
+ vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__a22o_1
X_14501_ net1410 vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11713_ net612 _07802_ _07907_ _07906_ vssd1 vssd1 vccd1 vccd1 _07908_ sky130_fd_sc_hd__a31o_2
XFILLER_0_16_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15481_ net1236 vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__inv_2
XANTENNA__12585__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12693_ net2567 net247 net385 vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17220_ clknet_leaf_82_wb_clk_i _02907_ _01203_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_14432_ net1227 vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_42_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11644_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\]
+ _07814_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] vssd1 vssd1 vccd1 vccd1
+ _07853_ sky130_fd_sc_hd__a31o_1
XFILLER_0_64_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17151_ clknet_leaf_43_wb_clk_i _02838_ _01134_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_3_5_0_wb_clk_i_X clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14363_ net1206 vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__inv_2
Xinput16 DAT_I[22] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10597__A0 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_30_Left_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11575_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[11\] _07784_ _07789_ vssd1 vssd1
+ vccd1 vccd1 _07792_ sky130_fd_sc_hd__and3_1
Xinput27 DAT_I[3] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16102_ clknet_leaf_138_wb_clk_i _01877_ _00090_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[9\]
+ sky130_fd_sc_hd__dfrtp_2
Xinput38 wb_rst_i vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_2
X_13314_ _07686_ _07708_ _03794_ net587 vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__o211a_1
X_17082_ clknet_leaf_76_wb_clk_i _02769_ _01065_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10526_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[31\] net676 net665 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06866_ sky130_fd_sc_hd__a22o_1
Xinput49 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__buf_1
X_14294_ net1346 vssd1 vssd1 vccd1 vccd1 _00088_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12338__A1 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13535__B1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16033_ clknet_leaf_139_wb_clk_i _01827_ _00027_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11929__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13245_ net2460 net355 net351 team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1
+ vccd1 vccd1 _01905_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10457_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[26\] net788 net751 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06797_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12889__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08370__Y _04710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09195__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09754__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13429__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13176_ net108 net848 net840 net1770 vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__a22o_1
X_10388_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[16\] net808 net774 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06728_ sky130_fd_sc_hd__a22o_1
XANTENNA__08530__C net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12127_ net2333 net218 net453 vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_5__f_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_5__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_17984_ net1499 vssd1 vssd1 vccd1 vccd1 la_data_out[26] sky130_fd_sc_hd__buf_2
XANTENNA__10134__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09923__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12058_ _07790_ net576 _07951_ vssd1 vssd1 vccd1 vccd1 _07955_ sky130_fd_sc_hd__and3_4
X_16935_ clknet_leaf_107_wb_clk_i _02622_ _00918_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11009_ _05707_ net512 vssd1 vssd1 vccd1 vccd1 _07349_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13445__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16866_ clknet_leaf_55_wb_clk_i _02553_ _00849_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_15817_ net1190 vssd1 vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16797_ clknet_leaf_70_wb_clk_i _02484_ _00780_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15748_ net1233 vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12813__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12495__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14015__B2 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15679_ net1317 vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__inv_2
XANTENNA__08493__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08220_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[61\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[53\]
+ net1051 vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__mux2_1
X_17418_ clknet_leaf_9_wb_clk_i _03105_ _01401_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11234__D1 _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08151_ net565 vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__inv_2
XANTENNA__08705__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17349_ clknet_leaf_47_wb_clk_i _03036_ _01332_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09442__A1 net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10309__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10052__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08082_ team_01_WB.instance_to_wrap.cpu.f0.i\[2\] _04555_ _04524_ vssd1 vssd1 vccd1
+ vccd1 _04556_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11839__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09745__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08984_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[8\] net670 _05321_ _05322_
+ _05323_ vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__a2111oi_1
XTAP_TAPCELL_ROW_149_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1017_A net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout477_A _07950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10331__X _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10512__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09605_ net996 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[24\] net971 vssd1
+ vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_27_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1386_A net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11068__A1 _05338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09536_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[28\] net790 net740 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09467_ _05760_ _05781_ net377 vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__o21ai_2
XANTENNA_fanout432_X net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout811_A net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout909_A _04785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08418_ net1026 net943 vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__nand2_4
XANTENNA__11603__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09398_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[27\] net698 net646 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08349_ net990 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[30\] net970 vssd1
+ vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__and3_1
XFILLER_0_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10043__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11360_ net1071 _07676_ _07682_ vssd1 vssd1 vccd1 vccd1 _07689_ sky130_fd_sc_hd__and3_1
XFILLER_0_61_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout899_X net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11749__S net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10311_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[18\] net811 net801 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06651_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11291_ _06886_ _06887_ _06960_ _04492_ vssd1 vssd1 vccd1 vccd1 _07631_ sky130_fd_sc_hd__a211o_1
XANTENNA__08631__B net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13030_ net2832 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[64\] net857 vssd1 vssd1
+ vccd1 vccd1 _02095_ sky130_fd_sc_hd__mux2_1
X_10242_ _06571_ _06579_ _06580_ _06581_ vssd1 vssd1 vccd1 vccd1 _06582_ sky130_fd_sc_hd__or4_1
XANTENNA__14190__B1 net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09446__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10173_ _06509_ _06510_ _06511_ _06512_ vssd1 vssd1 vccd1 vccd1 _06513_ sky130_fd_sc_hd__or4_1
XANTENNA__12721__X _03572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1103 net1115 vssd1 vssd1 vccd1 vccd1 net1103 sky130_fd_sc_hd__buf_2
Xfanout1114 net1115 vssd1 vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__buf_2
Xfanout1125 net1126 vssd1 vssd1 vccd1 vccd1 net1125 sky130_fd_sc_hd__clkbuf_2
Xfanout1136 net1141 vssd1 vssd1 vccd1 vccd1 net1136 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input38_A wb_rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1147 net1148 vssd1 vssd1 vccd1 vccd1 net1147 sky130_fd_sc_hd__clkbuf_2
X_14981_ net1254 vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__inv_2
XANTENNA__17733__Q team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout1158 net1160 vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__buf_2
XFILLER_0_156_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1169 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] vssd1 vssd1 vccd1 vccd1
+ net1169 sky130_fd_sc_hd__clkbuf_4
X_16720_ clknet_leaf_20_wb_clk_i _02407_ _00703_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout193 _07634_ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__buf_2
X_13932_ _04222_ _04223_ vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__nand2_2
XANTENNA__10503__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13863_ net1178 net1064 net2026 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[24\]
+ sky130_fd_sc_hd__and3b_1
X_16651_ clknet_leaf_9_wb_clk_i _02338_ _00634_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09181__C net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15602_ net1289 vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__inv_2
X_12814_ net1037 _07507_ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_83_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13794_ _04160_ _04162_ vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__nor2_1
X_16582_ clknet_leaf_90_wb_clk_i _02269_ _00565_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[14\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_69_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15533_ net1266 vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__inv_2
X_12745_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] net1060 net363 _03590_
+ vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10282__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15464_ net1375 vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__inv_2
X_12676_ net1972 net251 net390 vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14415_ net1342 vssd1 vssd1 vccd1 vccd1 _00209_ sky130_fd_sc_hd__inv_2
XANTENNA__08525__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17203_ clknet_leaf_23_wb_clk_i _02890_ _01186_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11627_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[26\] _07588_ net715 vssd1 vssd1
+ vccd1 vccd1 _07839_ sky130_fd_sc_hd__mux2_1
X_15395_ net1249 vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14346_ net1340 vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__inv_2
X_17134_ clknet_leaf_28_wb_clk_i _02821_ _01117_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11558_ net2880 _07786_ team_01_WB.instance_to_wrap.cpu.K0.count\[0\] vssd1 vssd1
+ vccd1 vccd1 _07788_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08822__A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold608 _01980_ vssd1 vssd1 vccd1 vccd1 net2143 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13508__B1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire583 _05865_ vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__buf_1
XFILLER_0_122_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17065_ clknet_leaf_36_wb_clk_i _02752_ _01048_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10509_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[31\] net734 _06831_ _06836_
+ _06839_ vssd1 vssd1 vccd1 vccd1 _06849_ sky130_fd_sc_hd__a2111o_1
Xhold619 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2154 sky130_fd_sc_hd__dlygate4sd3_1
X_14277_ net1343 vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__inv_2
X_11489_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[18\] net580 vssd1 vssd1 vccd1
+ vccd1 _07772_ sky130_fd_sc_hd__nand2_1
X_16016_ net1339 vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__inv_2
X_13228_ net2618 net352 net348 net1069 vssd1 vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__a22o_1
X_13159_ net1594 net847 _03734_ net1563 vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_55_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17967_ net1482 vssd1 vssd1 vccd1 vccd1 la_data_out[9] sky130_fd_sc_hd__buf_2
Xhold1308 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2843 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17643__Q team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold1319 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[23\] vssd1 vssd1 vccd1 vccd1
+ net2854 sky130_fd_sc_hd__dlygate4sd3_1
X_16918_ clknet_leaf_12_wb_clk_i _02605_ _00901_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_17898_ net1433 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_144_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09940__X _06280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_0_wb_clk_i sky130_fd_sc_hd__clkbuf_16
XANTENNA__09091__C net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16849_ clknet_leaf_114_wb_clk_i _02536_ _00832_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10030__C net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12798__A1 _07531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09321_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[24\] net657 net653 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[24\]
+ _05660_ vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__a221o_1
XANTENNA__13181__Y _03737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09252_ net1124 net711 net594 vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__a21o_1
X_08203_ net2840 net2723 net1042 vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09183_ net1009 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[16\] net883 vssd1
+ vssd1 vccd1 vccd1 _05523_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_32_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout225_A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08134_ _04600_ _04601_ _04602_ _04603_ vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__or4b_1
XANTENNA__11222__A1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10025__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09966__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08623__C1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13995__D _04286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08065_ _04538_ _04540_ _04541_ vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__or3_1
XANTENNA__08451__B net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1134_A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09718__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout594_A _04841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1301_A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10205__C net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09563__A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08967_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[8\] net665 _05304_ _05305_
+ _05306_ vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout761_A net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout382_X net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08898_ net1025 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[2\] net894 vssd1
+ vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout647_X net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10860_ _07198_ _07199_ net521 vssd1 vssd1 vccd1 vccd1 _07200_ sky130_fd_sc_hd__mux2_1
XANTENNA__08466__X _04806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08907__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12789__A1 _07553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13986__B1 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09519_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[29\] net798 net792 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout814_X net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10648__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10791_ _07100_ _07123_ _07124_ net327 _07130_ vssd1 vssd1 vccd1 vccd1 _07131_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12530_ net3074 net275 net404 vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__mux2_1
XANTENNA__11461__A1 net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_61_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12461_ net2331 net210 net411 vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__mux2_1
XANTENNA__12863__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13202__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14200_ _04154_ _04464_ vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__and2_1
XFILLER_0_136_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11412_ team_01_WB.instance_to_wrap.cpu.f0.i\[19\] _07692_ net323 vssd1 vssd1 vccd1
+ vccd1 _07729_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11213__A1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10016__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15180_ net1258 vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09738__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12392_ net2601 net221 net419 vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__mux2_1
XANTENNA__08642__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14131_ _04342_ _04396_ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_104_Left_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11343_ team_01_WB.instance_to_wrap.cpu.f0.i\[1\] _07671_ vssd1 vssd1 vccd1 vccd1
+ _07672_ sky130_fd_sc_hd__and2_1
XANTENNA__09709__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14062_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[83\] _04245_ _04247_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[67\]
+ _04350_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11274_ net557 _07498_ vssd1 vssd1 vccd1 vccd1 _07614_ sky130_fd_sc_hd__or2_1
XANTENNA__09176__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13013_ net3019 net3000 net865 vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__mux2_1
X_10225_ _05338_ _06564_ vssd1 vssd1 vccd1 vccd1 _06565_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_33_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09590__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09473__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17821_ clknet_leaf_95_wb_clk_i _03497_ _01761_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[91\]
+ sky130_fd_sc_hd__dfrtp_1
X_10156_ net340 vssd1 vssd1 vccd1 vccd1 _06496_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[25\] vssd1 vssd1 vccd1 vccd1 net1540
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12103__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17752_ clknet_leaf_116_wb_clk_i _03428_ _01692_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10087_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[7\] net741 _06413_ _06414_
+ _06415_ vssd1 vssd1 vccd1 vccd1 _06427_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10412__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14964_ net1379 vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_50_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16703_ clknet_leaf_43_wb_clk_i _02390_ _00686_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13915_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[7\] _04185_ _04204_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_113_Left_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17683_ clknet_leaf_129_wb_clk_i _03367_ _01624_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_14895_ net1388 vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload3_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14819__A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11942__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16634_ clknet_leaf_76_wb_clk_i _02321_ _00617_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13846_ net1180 net1066 net3176 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[7\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13442__B _05456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13977__B1 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13777_ _04162_ vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__inv_2
X_16565_ clknet_leaf_157_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[31\]
+ _00548_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10989_ _07005_ _07007_ vssd1 vssd1 vccd1 vccd1 _07329_ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15516_ net1246 vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12728_ _04510_ _03578_ vssd1 vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16496_ clknet_leaf_151_wb_clk_i _02250_ _00479_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12773__S net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12659_ net2576 net212 net387 vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__mux2_1
X_15447_ net1243 vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10007__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15378_ net1292 vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__inv_2
XANTENNA__17638__Q team_01_WB.instance_to_wrap.cpu.IG0.Instr\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12952__A1 _05300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17117_ clknet_leaf_64_wb_clk_i _02804_ _01100_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold405 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1940 sky130_fd_sc_hd__dlygate4sd3_1
X_14329_ net1202 vssd1 vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_57_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold416 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1951 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08620__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold427 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[13\] vssd1 vssd1 vccd1 vccd1
+ net1962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold438 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1973 sky130_fd_sc_hd__dlygate4sd3_1
X_17048_ clknet_leaf_61_wb_clk_i _02735_ _01031_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold449 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1984 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09086__C _04779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09870_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[12\] net805 net785 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06210_ sky130_fd_sc_hd__a22o_1
Xfanout907 net908 vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_74_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout918 _04775_ vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_146_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout929 net933 vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_146_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ net1024 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[1\] net933 vssd1
+ vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__and3_1
XFILLER_0_104_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1105 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[95\] vssd1 vssd1 vccd1 vccd1
+ net2640 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1116 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2651 sky130_fd_sc_hd__dlygate4sd3_1
X_08752_ net1012 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[4\] net910 vssd1
+ vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__and3_1
Xhold1127 _03465_ vssd1 vssd1 vccd1 vccd1 net2662 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1138 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2673 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10322__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12013__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1149 _01914_ vssd1 vssd1 vccd1 vccd1 net2684 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08136__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09333__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08683_ net1006 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[7\] net917 vssd1
+ vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__and3_1
XANTENNA__11140__A0 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11852__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14729__A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11691__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1084_A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09304_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[22\] net650 _05623_ _05624_
+ _05633_ vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10246__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11443__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_152_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10797__A3 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09235_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[21\] net663 net651 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__a22o_1
XANTENNA__12683__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout607_A _03583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout228_X net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1349_A net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09166_ net1010 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[16\] net900
+ vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__and3_1
XANTENNA__09939__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08462__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08117_ team_01_WB.instance_to_wrap.cpu.f0.i\[4\] team_01_WB.instance_to_wrap.cpu.f0.num\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__and2_1
XANTENNA__12943__A1 _05373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09097_ net1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[13\] net879
+ vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__and3_1
XANTENNA__10056__X _06396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_1__f_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1137_X net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14145__B1 _04258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08048_ net2063 net570 net346 net1072 vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold950 team_01_WB.instance_to_wrap.cpu.f0.num\[8\] vssd1 vssd1 vccd1 vccd1 net2485
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout597_X net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold961 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2496 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold972 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2507 sky130_fd_sc_hd__dlygate4sd3_1
Xhold983 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[22\] vssd1 vssd1 vccd1 vccd1
+ net2518 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1304_X net1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold994 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[57\] vssd1 vssd1 vccd1 vccd1
+ net2529 sky130_fd_sc_hd__dlygate4sd3_1
X_10010_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[1\] net800 net789 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06350_ sky130_fd_sc_hd__a22o_1
XANTENNA__09293__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09999_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] net626 _06337_ _06338_
+ vssd1 vssd1 vccd1 vccd1 _06339_ sky130_fd_sc_hd__a22o_2
XANTENNA_fanout764_X net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11636__A1_N net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1650 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 net3185
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09324__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11961_ net2390 net222 net471 vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__mux2_1
XANTENNA__12858__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout931_X net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13671__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11762__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13700_ team_01_WB.instance_to_wrap.cpu.c0.count\[9\] _04105_ vssd1 vssd1 vccd1 vccd1
+ _04121_ sky130_fd_sc_hd__or2_1
X_10912_ _06469_ _06472_ _06568_ _06566_ vssd1 vssd1 vccd1 vccd1 _07252_ sky130_fd_sc_hd__o31a_1
X_14680_ net1204 vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__inv_2
X_11892_ net575 _07942_ _07946_ vssd1 vssd1 vccd1 vccd1 _07949_ sky130_fd_sc_hd__and3_4
XANTENNA__08637__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13631_ _04051_ _04068_ vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_50_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10843_ _07139_ _07182_ net525 vssd1 vssd1 vccd1 vccd1 _07183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10237__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16350_ clknet_leaf_87_wb_clk_i _02104_ _00333_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[73\]
+ sky130_fd_sc_hd__dfrtp_1
X_13562_ _03921_ _03922_ vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__xor2_1
XFILLER_0_94_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10774_ _06712_ _06740_ _07112_ _06713_ _06677_ vssd1 vssd1 vccd1 vccd1 _07114_ sky130_fd_sc_hd__a311o_1
XANTENNA__11434__B2 _04483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12513_ net2089 net301 net408 vssd1 vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__mux2_1
X_15301_ net1286 vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__inv_2
X_16281_ clknet_leaf_125_wb_clk_i _02035_ _00264_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[4\]
+ sky130_fd_sc_hd__dfstp_1
X_13493_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[31\] _03953_ vssd1 vssd1
+ vccd1 vccd1 _03954_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12593__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08850__A2 _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15232_ net1233 vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__inv_2
X_12444_ net2948 net226 net415 vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08372__A team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08803__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12934__A1 _05415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15163_ net1253 vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__inv_2
X_12375_ net2157 net257 net426 vssd1 vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__mux2_1
XANTENNA__10945__A0 _06129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14114_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[70\] _04233_ _04236_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[54\]
+ _04399_ vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__a221o_1
XANTENNA__14136__B1 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11326_ _04548_ _07652_ _07660_ net1176 vssd1 vssd1 vccd1 vccd1 _07661_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15094_ net1261 vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__inv_2
XANTENNA__11937__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14045_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[91\] _04240_ _04243_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[27\]
+ _04333_ vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__a221o_1
X_11257_ _07592_ _07593_ _07595_ _07596_ vssd1 vssd1 vccd1 vccd1 _07597_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_52_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10208_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[8\] net821 _06535_ _06536_
+ _06544_ vssd1 vssd1 vccd1 vccd1 _06548_ sky130_fd_sc_hd__a2111o_1
X_11188_ _06979_ _07240_ vssd1 vssd1 vccd1 vccd1 _07528_ sky130_fd_sc_hd__nand2_1
XANTENNA__09634__C net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17804_ clknet_leaf_91_wb_clk_i net2360 _01744_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[74\]
+ sky130_fd_sc_hd__dfrtp_1
X_10139_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[11\] net799 net772 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06479_ sky130_fd_sc_hd__a22o_1
XANTENNA__08118__A1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13647__C1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15996_ net1368 vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_141_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17735_ clknet_leaf_116_wb_clk_i _03411_ _01675_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[5\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_141_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14947_ net1270 vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17666_ clknet_leaf_3_wb_clk_i _03351_ _01607_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_14878_ net1345 vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16617_ clknet_leaf_38_wb_clk_i _02304_ _00600_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16537__Q team_01_WB.instance_to_wrap.cpu.DM0.data_i\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13829_ net1660 net830 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[22\]
+ sky130_fd_sc_hd__and2_1
X_17597_ clknet_leaf_89_wb_clk_i _03284_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10859__S0 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16548_ clknet_leaf_1_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[14\]
+ _00531_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16479_ clknet_leaf_151_wb_clk_i _02233_ _00462_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08841__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09020_ net1095 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[9\] net910 vssd1
+ vssd1 vccd1 vccd1 _05360_ sky130_fd_sc_hd__and3_1
XANTENNA__11260__X _07600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11189__B1 _07528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12925__A1 _03692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08713__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12008__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold202 team_01_WB.instance_to_wrap.cpu.f0.write_data\[21\] vssd1 vssd1 vccd1 vccd1
+ net1737 sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[107\] vssd1 vssd1 vccd1 vccd1
+ net1748 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14127__B1 _04254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold224 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[127\] vssd1 vssd1 vccd1 vccd1
+ net1759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[0\] vssd1 vssd1 vccd1 vccd1 net1770
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1781 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold257 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1792 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 _02014_ vssd1 vssd1 vccd1 vccd1 net1803 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11847__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09922_ net1153 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[4\] net974 vssd1
+ vssd1 vccd1 vccd1 _06262_ sky130_fd_sc_hd__and3_1
XANTENNA__12091__X _07956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold279 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1814 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout704 _04758_ vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__buf_4
Xfanout715 net717 vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__clkbuf_4
Xfanout726 net728 vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09554__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout737 net738 vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__buf_6
X_09853_ net373 _06191_ vssd1 vssd1 vccd1 vccd1 _06193_ sky130_fd_sc_hd__nand2_1
Xfanout748 _04682_ vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__buf_4
Xfanout759 net762 vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__clkbuf_8
X_08804_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[0\] net674 _05141_ _05142_
+ _05143_ vssd1 vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__a2111o_1
X_09784_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[15\] _04634_ net800
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[15\] vssd1 vssd1 vccd1 vccd1
+ _06124_ sky130_fd_sc_hd__a22o_1
XANTENNA__13638__C1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08735_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\] net599 net596 vssd1 vssd1
+ vccd1 vccd1 _05075_ sky130_fd_sc_hd__and3_1
XANTENNA__12678__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout557_A net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1299_A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08666_ _04971_ _05005_ net602 vssd1 vssd1 vccd1 vccd1 _05006_ sky130_fd_sc_hd__mux2_2
XANTENNA__10467__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08597_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[15\] net943 net663 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[15\]
+ net706 vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout724_A net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1087_X net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10219__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_134_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_48_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout512_X net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08463__Y _04803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09490__C1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_779 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09218_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[17\] net676 _05531_
+ _05539_ _05540_ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10490_ net1130 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[31\] net951
+ vssd1 vssd1 vccd1 vccd1 _06830_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_20_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12916__A1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09149_ _05480_ _05481_ _05487_ _05488_ vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__or4_1
XFILLER_0_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10927__B1 _07265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10227__A _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14118__B1 _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12160_ net2255 net219 net449 vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout881_X net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11111_ _06404_ _06405_ _07450_ vssd1 vssd1 vccd1 vccd1 _07451_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout979_X net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10942__A3 _06738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12091_ _07791_ net575 _07945_ vssd1 vssd1 vccd1 vccd1 _07956_ sky130_fd_sc_hd__and3_4
Xhold780 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2315 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold791 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2326 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09545__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11042_ _05076_ _06250_ vssd1 vssd1 vccd1 vccd1 _07382_ sky130_fd_sc_hd__nor2_1
XANTENNA__10155__A1 _06494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15850_ net1334 vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14801_ net1395 vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__inv_2
XANTENNA_input20_A DAT_I[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15781_ net1203 vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__inv_2
XANTENNA__09848__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13644__A2 _07323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12993_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[93\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[101\]
+ net860 vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__mux2_1
X_17520_ clknet_leaf_146_wb_clk_i _03207_ _01503_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1480 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[19\] vssd1 vssd1 vccd1 vccd1
+ net3015 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11655__A1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14732_ net1210 vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__inv_2
Xhold1491 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[32\] vssd1 vssd1 vccd1 vccd1
+ net3026 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11944_ net1856 net253 net476 vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__mux2_1
XANTENNA__08367__A _04706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11505__B _07756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17451_ clknet_leaf_7_wb_clk_i _03138_ _01434_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11875_ net2127 net262 net484 vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__mux2_1
X_14663_ net1305 vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16402_ clknet_leaf_100_wb_clk_i _02156_ _00385_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[125\]
+ sky130_fd_sc_hd__dfstp_1
X_10826_ net333 net336 _07164_ vssd1 vssd1 vccd1 vccd1 _07166_ sky130_fd_sc_hd__mux2_1
X_13614_ _03887_ _04054_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__xnor2_1
X_17382_ clknet_leaf_90_wb_clk_i _03069_ _01365_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14594_ net1358 vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_45_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16333_ clknet_leaf_122_wb_clk_i _02087_ _00316_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[56\]
+ sky130_fd_sc_hd__dfrtp_1
X_10757_ _04844_ net510 net333 _07096_ vssd1 vssd1 vccd1 vccd1 _07097_ sky130_fd_sc_hd__a31o_1
X_13545_ _03928_ _03991_ vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17899__1434 vssd1 vssd1 vccd1 vccd1 _17899__1434/HI net1434 sky130_fd_sc_hd__conb_1
XANTENNA__10091__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09198__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13476_ _04500_ _04842_ _03927_ vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__o21ba_1
X_16264_ clknet_leaf_141_wb_clk_i net1718 _00252_ vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10688_ _06891_ _06937_ net533 vssd1 vssd1 vccd1 vccd1 _07028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09629__C net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18003_ net1507 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__buf_2
XANTENNA__12907__A1 _05615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15215_ net1386 vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__inv_2
X_12427_ net2374 net216 net417 vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16195_ clknet_leaf_159_wb_clk_i _01955_ _00183_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12904__X _03678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14832__A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13580__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09784__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12358_ net2796 net188 net423 vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__mux2_1
X_15146_ net1374 vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__inv_2
XANTENNA__08830__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11667__S net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11309_ net727 _07438_ _07647_ vssd1 vssd1 vccd1 vccd1 _07648_ sky130_fd_sc_hd__a21o_1
X_15077_ net1262 vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_71_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12289_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[1\] net314 net437 vssd1
+ vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14028_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[106\] _04252_ _04315_ _04317_
+ vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__a211o_1
XANTENNA__09536__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13332__B2 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11239__Y _07579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_0__f_wb_clk_i_X clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_101_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12498__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15979_ net1413 vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__inv_2
XANTENNA__13635__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13183__A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08520_ net1081 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[18\] net897
+ vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__and3_1
X_17718_ clknet_leaf_115_wb_clk_i _03402_ _01659_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08451_ net1108 net944 vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__and2_2
XANTENNA__08708__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17649_ clknet_leaf_15_wb_clk_i _03334_ _01590_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08382_ net1170 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[4\]
+ _04711_ vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__nor4_1
XFILLER_0_129_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09067__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14060__A2 _04236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08814__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_118_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_118_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_143_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10621__A2 _06887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09539__C net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09003_ net1094 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[9\] net887 vssd1
+ vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11150__B _07489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout305_A _07935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13571__A1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09775__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08740__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout501 net502 vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__buf_6
XANTENNA__09527__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09905_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[5\] net822 net796 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06245_ sky130_fd_sc_hd__a22o_1
Xfanout512 _05931_ vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__buf_4
XFILLER_0_10_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout523 net526 vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__buf_2
Xfanout534 _05190_ vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout674_A _04791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout295_X net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout545 _05152_ vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__clkbuf_2
Xfanout556 _05114_ vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__clkbuf_4
X_09836_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[13\] net755 net754 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06176_ sky130_fd_sc_hd__a22o_1
Xfanout567 net568 vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__buf_2
Xfanout578 _07753_ vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1002_X net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout589 _07785_ vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13087__A0 _03710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout462_X net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09767_ _06002_ _06036_ _06104_ _06106_ vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout841_A net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout939_A net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08718_ net1097 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[5\] net941 vssd1
+ vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__and3_1
XANTENNA__12201__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09698_ net996 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[21\] net979 vssd1
+ vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08502__A1 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08649_ net1020 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[10\] net912
+ vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout727_X net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11660_ net611 _07815_ _07865_ _07864_ vssd1 vssd1 vccd1 vccd1 _07866_ sky130_fd_sc_hd__a31o_2
XTAP_TAPCELL_ROW_25_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14051__A2 _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10611_ net546 _06313_ vssd1 vssd1 vccd1 vccd1 _06951_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11591_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\]
+ _07805_ vssd1 vssd1 vccd1 vccd1 _07808_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13330_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[18\] net826 _03806_ _03807_
+ vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__o22a_1
X_10542_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] _06881_ net600 vssd1 vssd1
+ vccd1 vccd1 _06882_ sky130_fd_sc_hd__mux2_4
XFILLER_0_135_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13261_ _04470_ _03752_ vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_40_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10473_ _05729_ _05736_ vssd1 vssd1 vccd1 vccd1 _06813_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_40_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12212_ net2560 net252 net446 vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__mux2_1
X_15000_ net1213 vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13192_ net17 net835 net628 net2241 vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__o22a_1
XANTENNA__08650__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input68_A wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12143_ net2355 net254 net452 vssd1 vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__mux2_1
XANTENNA__13268__A team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10915__A3 _06158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_4__f_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_4__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09518__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12074_ net2181 net264 net461 vssd1 vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__mux2_1
X_16951_ clknet_leaf_14_wb_clk_i _02638_ _00934_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09184__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15902_ net1408 vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__inv_2
XANTENNA__15483__A net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11025_ _04948_ net374 vssd1 vssd1 vccd1 vccd1 _07365_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12900__A _05654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16882_ clknet_leaf_110_wb_clk_i _02569_ _00865_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10898__Y _07238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15833_ net1331 vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__inv_2
XANTENNA__13617__A2 _07207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08368__Y _04708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12111__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15764_ net1198 vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__inv_2
XANTENNA__10420__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12976_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[110\] net2960 net855 vssd1 vssd1
+ vccd1 vccd1 _02149_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17503_ clknet_leaf_43_wb_clk_i _03190_ _01486_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14715_ net1186 vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__inv_2
XANTENNA__08528__C net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11927_ net2811 net221 net475 vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__mux2_1
X_15695_ net1299 vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11950__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17434_ clknet_leaf_76_wb_clk_i _03121_ _01417_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14646_ net1231 vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__inv_2
X_11858_ net1843 net290 net487 vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14042__A2 _04265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08825__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_19 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_6_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10809_ net522 net518 vssd1 vssd1 vccd1 vccd1 _07149_ sky130_fd_sc_hd__nor2_1
X_17365_ clknet_leaf_111_wb_clk_i _03052_ _01348_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11789_ net1901 net316 net496 vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__mux2_1
XANTENNA__13843__A_N net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14577_ net1413 vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11251__A net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16316_ clknet_leaf_120_wb_clk_i _02070_ _00299_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13528_ net198 net194 _07846_ net644 vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_60_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17296_ clknet_leaf_147_wb_clk_i _02983_ _01279_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18011__1510 vssd1 vssd1 vccd1 vccd1 _18011__1510/HI net1510 sky130_fd_sc_hd__conb_1
XFILLER_0_125_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16247_ clknet_leaf_151_wb_clk_i net1640 _00235_ vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13459_ _03858_ _03919_ vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13553__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09757__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__buf_2
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__buf_2
X_16178_ clknet_leaf_1_wb_clk_i _01938_ _00166_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput126 net126 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__buf_2
XANTENNA__10367__B2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput137 net137 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__buf_2
XFILLER_0_140_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15129_ net1235 vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__inv_2
Xoutput148 net148 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
Xoutput159 net159 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
XANTENNA__10154__X _06494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09094__C net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09391__A net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09621_ _05952_ _05953_ _05957_ _05960_ vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_108_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13608__A2 _07520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09552_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[28\] net812 net749 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__a22o_1
XANTENNA__12021__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08503_ net1118 net711 net600 _04841_ vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__a211o_1
XFILLER_0_78_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09483_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[30\] net680 _05809_
+ _05811_ _05814_ vssd1 vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12956__S net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout255_A net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12809__X _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12831__A3 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11713__X _07908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11860__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08434_ net1082 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[23\] net922
+ vssd1 vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__and3_1
XANTENNA__08294__X _04634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14033__A2 _04245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08735__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13360__B net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08365_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[30\] net763 net623 vssd1
+ vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10329__X _06669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08454__B net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1164_A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08296_ net1153 net977 vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__and2_2
XANTENNA__09460__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12691__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1331_A net1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1429_A net1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13544__A1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout791_A net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08901__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout889_A net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_86_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout1307 net1310 vssd1 vssd1 vccd1 vccd1 net1307 sky130_fd_sc_hd__buf_4
Xfanout320 _07937_ vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_15_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout1318 net1321 vssd1 vssd1 vccd1 vccd1 net1318 sky130_fd_sc_hd__buf_4
XANTENNA_fanout677_X net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout331 _06923_ vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__clkbuf_4
Xfanout1329 net1332 vssd1 vssd1 vccd1 vccd1 net1329 sky130_fd_sc_hd__clkbuf_4
Xfanout353 _03741_ vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__buf_2
Xfanout364 _03580_ vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__clkbuf_4
Xfanout375 _05262_ vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__clkbuf_4
X_17898__1433 vssd1 vssd1 vccd1 vccd1 _17898__1433/HI net1433 sky130_fd_sc_hd__conb_1
XANTENNA__09920__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout386 _03570_ vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__clkbuf_4
X_09819_ _06158_ vssd1 vssd1 vccd1 vccd1 _06159_ sky130_fd_sc_hd__inv_2
Xfanout397 _03567_ vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__buf_6
XANTENNA__09732__C net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout844_X net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12830_ net1746 net641 net609 _03649_ vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11055__B _06280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12761_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[22\] _07154_ net1032 vssd1 vssd1
+ vccd1 vccd1 _03602_ sky130_fd_sc_hd__mux2_1
XANTENNA__13866__A_N net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11770__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14500_ net1406 vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11712_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] _07801_ vssd1 vssd1 vccd1
+ vccd1 _07907_ sky130_fd_sc_hd__or2_1
X_15480_ net1213 vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__inv_2
X_12692_ net2729 net213 net383 vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__mux2_1
XANTENNA__08645__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14024__A2 _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12035__A1 _07858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11643_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[23\] _07111_ net713 vssd1 vssd1
+ vccd1 vccd1 _07852_ sky130_fd_sc_hd__mux2_1
X_14431_ net1335 vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_42_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09436__C1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09987__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17150_ clknet_leaf_85_wb_clk_i _02837_ _01133_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14362_ net1336 vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__inv_2
X_11574_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\] team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\]
+ vssd1 vssd1 vccd1 vccd1 _07791_ sky130_fd_sc_hd__nor2_2
XANTENNA__09179__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10597__A1 _06158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput17 DAT_I[23] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09451__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16101_ clknet_leaf_127_wb_clk_i _01876_ _00089_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[8\]
+ sky130_fd_sc_hd__dfrtp_2
Xinput28 DAT_I[4] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
X_13313_ team_01_WB.instance_to_wrap.cpu.f0.i\[18\] net610 _07705_ team_01_WB.instance_to_wrap.cpu.f0.i\[19\]
+ vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__a31o_1
Xinput39 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
X_10525_ _06859_ _06860_ _06864_ vssd1 vssd1 vccd1 vccd1 _06865_ sky130_fd_sc_hd__or3_1
X_14293_ net1346 vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__inv_2
X_17081_ clknet_leaf_71_wb_clk_i _02768_ _01064_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13535__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13244_ net3136 net354 net350 team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1
+ vccd1 vccd1 _01906_ sky130_fd_sc_hd__a22o_1
X_16032_ clknet_leaf_131_wb_clk_i _01826_ net1185 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10456_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[26\] net740 _06783_ _06784_
+ _06785_ vssd1 vssd1 vccd1 vccd1 _06796_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_150_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11546__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13175_ net119 net848 net840 net2101 vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__a22o_1
XANTENNA__12106__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10387_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[16\] net801 net756 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06727_ sky130_fd_sc_hd__a22o_1
XANTENNA__10415__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12126_ net2577 net223 net451 vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__mux2_1
X_17983_ net1498 vssd1 vssd1 vccd1 vccd1 la_data_out[25] sky130_fd_sc_hd__buf_2
XANTENNA__11945__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16934_ clknet_leaf_72_wb_clk_i _02621_ _00917_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12057_ net2229 net288 net464 vssd1 vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__mux2_1
XANTENNA__10702__X _07042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11008_ _05707_ _05932_ vssd1 vssd1 vccd1 vccd1 _07348_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_88_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16865_ clknet_leaf_54_wb_clk_i _02552_ _00848_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_15816_ net1192 vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__inv_2
X_16796_ clknet_leaf_59_wb_clk_i _02483_ _00779_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15747_ net1251 vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__inv_2
X_12959_ net1874 net870 net357 _03714_ vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10285__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15678_ net1317 vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__inv_2
XANTENNA__14015__A2 _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17417_ clknet_leaf_40_wb_clk_i _03104_ _01400_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14629_ net1385 vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08150_ _04604_ _04619_ team_01_WB.instance_to_wrap.cpu.f0.state\[6\] _04516_ vssd1
+ vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__o211a_1
X_17348_ clknet_leaf_82_wb_clk_i _03035_ _01331_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09938__X _06278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09089__C net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_151_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08081_ _04531_ _04540_ _04545_ _04554_ vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__or4b_1
XANTENNA__15388__A net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17279_ clknet_leaf_41_wb_clk_i _02966_ _01262_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap1182 _07786_ vssd1 vssd1 vccd1 vccd1 net1182 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_3_0_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__16280__Q team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12016__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10325__A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08983_ net1088 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[8\] net929 vssd1
+ vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11855__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11708__X _07904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08289__X _04629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09902__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08449__B net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11156__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09604_ net1146 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[24\] net946
+ vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_27_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11068__A2 _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09535_ net996 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[28\] net985 vssd1
+ vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__and3_1
XANTENNA__12686__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1281_A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout637_A net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_133_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_133_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1379_A net1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09466_ _05805_ vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__inv_2
XANTENNA__14006__A2 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08465__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09681__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08417_ net1026 net943 vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09397_ _05659_ _05681_ _05707_ _05729_ net560 vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__a41o_1
XANTENNA__13214__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout804_A _04643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout425_X net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_502 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08348_ net991 net970 vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09848__X _06188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09433__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08279_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[2\] net1817 net1043 vssd1 vssd1
+ vccd1 vccd1 _03408_ sky130_fd_sc_hd__mux2_1
XANTENNA__13517__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10310_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[18\] net804 _06647_
+ _06648_ _06649_ vssd1 vssd1 vccd1 vccd1 _06650_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_21_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09296__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11290_ net1169 _04712_ vssd1 vssd1 vccd1 vccd1 _07630_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout794_X net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10241_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[9\] net813 net732 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06581_ sky130_fd_sc_hd__a22o_1
X_10172_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[10\] _04636_ net810
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[10\] vssd1 vssd1 vccd1 vccd1
+ _06512_ sky130_fd_sc_hd__a22o_1
Xfanout1104 net1106 vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__buf_2
Xfanout1115 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[24\] vssd1 vssd1 vccd1 vccd1
+ net1115 sky130_fd_sc_hd__buf_4
XANTENNA__11765__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1126 net1127 vssd1 vssd1 vccd1 vccd1 net1126 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1137 net1141 vssd1 vssd1 vccd1 vccd1 net1137 sky130_fd_sc_hd__buf_2
X_14980_ net1233 vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_35_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1148 net1151 vssd1 vssd1 vccd1 vccd1 net1148 sky130_fd_sc_hd__clkbuf_2
Xfanout1159 net1160 vssd1 vssd1 vccd1 vccd1 net1159 sky130_fd_sc_hd__buf_1
X_13931_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[3\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__and2b_2
Xfanout194 _07634_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__clkbuf_4
X_16650_ clknet_leaf_32_wb_clk_i _02337_ _00633_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13862_ net1177 net1064 net2789 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[23\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_69_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15601_ net1394 vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__inv_2
X_12813_ net1828 net640 net608 _03637_ vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_2_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16581_ clknet_leaf_50_wb_clk_i _02268_ _00564_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_2_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12596__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13793_ _04156_ _01833_ vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15532_ net1259 vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12744_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[27\] _07566_ net1034 vssd1 vssd1
+ vccd1 vccd1 _03590_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08806__C net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15463_ net1389 vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13205__B1 _03738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12675_ net3039 net226 net387 vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__mux2_1
XANTENNA__10019__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17202_ clknet_leaf_110_wb_clk_i _02889_ _01185_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14414_ net1323 vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__inv_2
XANTENNA__09758__X _06098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11626_ net3116 net213 net499 vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__mux2_1
X_15394_ net1321 vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__inv_2
XANTENNA__09424__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17133_ clknet_leaf_108_wb_clk_i _02820_ _01116_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14345_ net1330 vssd1 vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__inv_2
X_11557_ net2778 _07787_ vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__xor2_1
XFILLER_0_107_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold609 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2144 sky130_fd_sc_hd__dlygate4sd3_1
Xwire584 _05453_ vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__clkbuf_4
X_17064_ clknet_leaf_62_wb_clk_i _02751_ _01047_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10508_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[31\] net776 net752 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[31\]
+ _06843_ vssd1 vssd1 vccd1 vccd1 _06848_ sky130_fd_sc_hd__a221o_1
XFILLER_0_80_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11488_ net367 _07771_ net3010 net875 vssd1 vssd1 vccd1 vccd1 _03350_ sky130_fd_sc_hd__o2bb2a_1
X_14276_ net1340 vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__inv_2
XANTENNA__09637__C net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16015_ net1341 vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_59_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10439_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] net627 _06777_ _06778_
+ vssd1 vssd1 vccd1 vccd1 _06779_ sky130_fd_sc_hd__a22o_2
X_13227_ net2947 net353 net349 team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1
+ vccd1 vccd1 _01923_ sky130_fd_sc_hd__a22o_1
X_17928__1535 vssd1 vssd1 vccd1 vccd1 net1535 _17928__1535/LO sky130_fd_sc_hd__conb_1
X_13158_ net1595 net846 net839 net1557 vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_55_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11675__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12109_ net2431 net258 net457 vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__mux2_1
X_17966_ net1481 vssd1 vssd1 vccd1 vccd1 la_data_out[8] sky130_fd_sc_hd__buf_2
X_13089_ _03712_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[5\] net853 vssd1 vssd1
+ vccd1 vccd1 _02036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1309 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2844 sky130_fd_sc_hd__dlygate4sd3_1
X_16917_ clknet_leaf_118_wb_clk_i _02604_ _00900_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_17897_ net1432 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_144_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16848_ clknet_leaf_144_wb_clk_i _02535_ _00831_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16779_ clknet_leaf_9_wb_clk_i _02466_ _00762_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09320_ net1115 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[24\] net909
+ net647 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[24\] vssd1 vssd1 vccd1
+ vccd1 _05660_ sky130_fd_sc_hd__a32o_1
XFILLER_0_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08716__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09251_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[21\] net703 _05585_ _05590_
+ vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__o22a_4
XANTENNA__08871__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08202_ net2756 net2712 net1048 vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__mux2_1
XANTENNA__13747__A1 _04504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09182_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[16\] net658 _05519_
+ _05520_ _05521_ vssd1 vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_7_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08133_ _04477_ team_01_WB.instance_to_wrap.cpu.f0.num\[17\] team_01_WB.instance_to_wrap.cpu.f0.num\[6\]
+ _04487_ _04594_ vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_32_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17897__1432 vssd1 vssd1 vccd1 vccd1 _17897__1432/HI net1432 sky130_fd_sc_hd__conb_1
XFILLER_0_114_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout218_A _07831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08064_ _04514_ _04529_ vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_79_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08966_ net1087 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[8\] net911 vssd1
+ vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__and3_1
XANTENNA__09282__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08897_ net1025 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[2\] net890 vssd1
+ vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout375_X net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10497__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_40_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout542_X net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09518_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[29\] net802 net731 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[29\]
+ _05846_ vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__a221o_1
XFILLER_0_151_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10790_ net515 _06957_ _07099_ _07129_ vssd1 vssd1 vccd1 vccd1 _07130_ sky130_fd_sc_hd__a31o_1
XFILLER_0_13_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09449_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[29\] net700 net655 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout807_X net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12460_ net2813 net215 net413 vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__mux2_1
XANTENNA__09406__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11411_ _07701_ _07709_ _07728_ net323 vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12391_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[31\] net191 net419 vssd1
+ vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__mux2_1
XANTENNA__08614__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10517__X _06857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11342_ team_01_WB.instance_to_wrap.cpu.f0.i\[0\] net1175 _07670_ vssd1 vssd1 vccd1
+ vccd1 _07671_ sky130_fd_sc_hd__and3_1
X_14130_ net1756 net604 _04415_ net1185 vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_30_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11273_ _06100_ _07089_ _06104_ vssd1 vssd1 vccd1 vccd1 _07613_ sky130_fd_sc_hd__a21o_1
X_14061_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[43\] _04246_ _04264_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[107\]
+ vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13012_ net2802 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[82\] net863 vssd1 vssd1
+ vccd1 vccd1 _02113_ sky130_fd_sc_hd__mux2_1
XANTENNA_input50_A wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10224_ _05264_ _05265_ _05302_ _04750_ vssd1 vssd1 vccd1 vccd1 _06564_ sky130_fd_sc_hd__o31a_1
X_17820_ clknet_leaf_91_wb_clk_i _03496_ _01760_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[90\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_33_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10155_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] _06494_ net623 vssd1
+ vssd1 vccd1 vccd1 _06495_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_33_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16530__CLK clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17751_ clknet_leaf_98_wb_clk_i _03427_ _01691_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[21\]
+ sky130_fd_sc_hd__dfstp_1
X_10086_ _06422_ _06423_ _06424_ _06425_ vssd1 vssd1 vccd1 vccd1 _06426_ sky130_fd_sc_hd__or4_1
X_14963_ net1392 vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__inv_2
XANTENNA__09192__C net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold6 team_01_WB.instance_to_wrap.cpu.f0.write_data\[0\] vssd1 vssd1 vccd1 vccd1
+ net1541 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12477__A1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16702_ clknet_leaf_80_wb_clk_i _02389_ _00685_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13914_ net2875 _04209_ _04210_ vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__o21a_1
X_17682_ clknet_leaf_129_wb_clk_i _03366_ _01623_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_89_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14894_ net1297 vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_18_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16633_ clknet_leaf_102_wb_clk_i _02320_ _00616_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13845_ net1179 net1066 net1601 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[6\]
+ sky130_fd_sc_hd__and3b_1
X_16564_ clknet_leaf_158_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[30\]
+ _00547_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13776_ net1184 _04161_ vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__nand2_2
XFILLER_0_57_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10988_ net540 _07327_ vssd1 vssd1 vccd1 vccd1 _07328_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09645__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15515_ net1275 vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__inv_2
X_12727_ net1033 _03576_ _03577_ net1175 vssd1 vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__a211o_1
XFILLER_0_127_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16495_ clknet_leaf_141_wb_clk_i _02249_ _00478_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12907__X _03680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15446_ net1261 vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12658_ net2887 net216 net389 vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11609_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] _07820_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\]
+ vssd1 vssd1 vccd1 vccd1 _07825_ sky130_fd_sc_hd__a21o_1
X_15377_ net1393 vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12589_ net2159 net190 net395 vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17116_ clknet_leaf_59_wb_clk_i _02803_ _01099_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14328_ net1189 vssd1 vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_57_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold406 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1941 sky130_fd_sc_hd__dlygate4sd3_1
Xhold417 net135 vssd1 vssd1 vccd1 vccd1 net1952 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold428 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1963 sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[8\] vssd1 vssd1 vccd1 vccd1 net1974
+ sky130_fd_sc_hd__dlygate4sd3_1
X_17047_ clknet_leaf_13_wb_clk_i _02734_ _01030_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14259_ net1205 vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09664__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout908 net909 vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__clkbuf_4
Xfanout919 net920 vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[1\] net692 net675 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_146_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1106 _03501_ vssd1 vssd1 vccd1 vccd1 net2641 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1117 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2652 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2663 sky130_fd_sc_hd__dlygate4sd3_1
X_08751_ net1099 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[4\] net921 vssd1
+ vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__and3_1
XFILLER_0_139_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17949_ net1464 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
Xhold1139 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2674 sky130_fd_sc_hd__dlygate4sd3_1
X_08682_ net1086 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[7\] net896 vssd1
+ vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__and3_1
XANTENNA__11140__A1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10041__C net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14090__B1 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09303_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[22\] net935
+ vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__and3_1
XANTENNA__08446__C net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11443__A2 team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12964__S net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_124_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout335_A _06912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1077_A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09234_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[21\] net697 net647 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08743__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09165_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[16\] net693 net667 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[16\]
+ _05504_ vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13196__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1244_A net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08116_ team_01_WB.instance_to_wrap.cpu.f0.i\[4\] team_01_WB.instance_to_wrap.cpu.f0.num\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12943__A2 _07757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09096_ net1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[13\] net896
+ vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__and3_1
XANTENNA__11600__C team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08611__A3 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08047_ net1669 net569 net347 net1070 vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1032_X net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold940 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold951 _01908_ vssd1 vssd1 vccd1 vccd1 net2486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold973 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2508 sky130_fd_sc_hd__dlygate4sd3_1
Xhold984 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2519 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout492_X net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout871_A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold995 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2530 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout969_A _04648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12204__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10182__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[2\] net765 net624 vssd1
+ vssd1 vccd1 vccd1 _06338_ sky130_fd_sc_hd__o21a_1
XANTENNA__09309__D1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12459__A1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08949_ net1027 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[6\] net937 vssd1
+ vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_4_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout757_X net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13120__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1640 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 net3175
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1651 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[14\] vssd1 vssd1 vccd1 vccd1
+ net3186 sky130_fd_sc_hd__dlygate4sd3_1
X_11960_ net2922 net189 net471 vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__mux2_1
XANTENNA__08477__X _04817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10911_ _07114_ _07233_ _07239_ _07250_ vssd1 vssd1 vccd1 vccd1 _07251_ sky130_fd_sc_hd__a211o_2
X_11891_ net1790 net288 net483 vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout924_X net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09740__C net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11344__A team_01_WB.instance_to_wrap.cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13630_ _03883_ _03895_ vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__nand2_1
X_10842_ _07180_ _07181_ net520 vssd1 vssd1 vccd1 vccd1 _07182_ sky130_fd_sc_hd__mux2_1
XANTENNA__14081__B1 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12631__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13561_ net986 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] _04009_ _04010_
+ vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__a22o_1
XANTENNA__08835__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10773_ _06712_ _06740_ _07112_ _06713_ vssd1 vssd1 vccd1 vccd1 _07113_ sky130_fd_sc_hd__a31o_1
X_17927__1534 vssd1 vssd1 vccd1 vccd1 net1534 _17927__1534/LO sky130_fd_sc_hd__conb_1
XFILLER_0_94_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10642__A0 _06129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15300_ net1230 vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__inv_2
X_12512_ net2128 net282 net410 vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__mux2_1
X_16280_ clknet_leaf_125_wb_clk_i _02034_ _00263_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08653__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13492_ net710 _04729_ net596 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1
+ vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__o31a_1
XANTENNA__13187__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15231_ net1312 vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12443_ net3003 net284 net418 vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08372__B team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12934__A2 _07757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15162_ net1371 vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09260__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12374_ net2688 net230 net425 vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__mux2_1
XANTENNA__10945__A1 _06158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14113_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[6\] _04265_ _04266_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__a22o_1
X_11325_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[4\] _07659_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[5\]
+ vssd1 vssd1 vccd1 vccd1 _07660_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_95_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15093_ net1275 vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11256_ _05681_ net330 _07350_ net368 _07591_ vssd1 vssd1 vccd1 vccd1 _07596_ sky130_fd_sc_hd__o221a_1
X_14044_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[83\] _04251_ _04266_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08366__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10207_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[8\] net779 net739 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _06547_ sky130_fd_sc_hd__a22o_1
XANTENNA__12114__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11187_ net530 _07237_ vssd1 vssd1 vccd1 vccd1 _07527_ sky130_fd_sc_hd__or2_1
X_17803_ clknet_leaf_94_wb_clk_i net2676 _01743_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[73\]
+ sky130_fd_sc_hd__dfrtp_1
X_10138_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[11\] net759 _06476_
+ _06477_ vssd1 vssd1 vccd1 vccd1 _06478_ sky130_fd_sc_hd__a211o_1
X_15995_ net1364 vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__inv_2
XANTENNA__11953__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09315__A1 net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17734_ clknet_leaf_116_wb_clk_i _03410_ _01674_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[4\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_141_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10069_ _06406_ _06408_ vssd1 vssd1 vccd1 vccd1 _06409_ sky130_fd_sc_hd__nor2_1
X_14946_ net1320 vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_141_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17896__1431 vssd1 vssd1 vccd1 vccd1 _17896__1431/HI net1431 sky130_fd_sc_hd__conb_1
XANTENNA__11122__A1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09866__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11122__B2 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17665_ clknet_leaf_0_wb_clk_i _03350_ _01606_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14877_ net1240 vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__inv_2
X_16616_ clknet_leaf_61_wb_clk_i _02303_ _00599_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13828_ net3006 net831 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[21\]
+ sky130_fd_sc_hd__and2_1
X_17596_ clknet_leaf_86_wb_clk_i _03283_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09618__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14072__B1 _04266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16547_ clknet_leaf_2_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[13\]
+ _00530_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13759_ _04147_ vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_139_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09659__A net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16478_ clknet_leaf_151_wb_clk_i _02232_ _00461_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08563__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15429_ net1255 vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__inv_2
XANTENNA__13178__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16576__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08850__X _05190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09097__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold203 team_01_WB.instance_to_wrap.a1.ADR_I\[13\] vssd1 vssd1 vccd1 vccd1 net1738
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 _03521_ vssd1 vssd1 vccd1 vccd1 net1749 sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 _03533_ vssd1 vssd1 vccd1 vccd1 net1760 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold236 _01966_ vssd1 vssd1 vccd1 vccd1 net1771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[123\] vssd1 vssd1 vccd1 vccd1
+ net1782 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10036__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold258 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1793 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[4\] net804 net733 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06261_ sky130_fd_sc_hd__a22o_1
XANTENNA__09394__A net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold269 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1804 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout705 net708 vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08357__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout716 net717 vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12024__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09852_ net373 _06191_ vssd1 vssd1 vccd1 vccd1 _06192_ sky130_fd_sc_hd__nor2_1
Xfanout727 net728 vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__clkbuf_4
Xfanout738 _04686_ vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__buf_6
XANTENNA__10333__A net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout749 _04680_ vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__buf_6
XFILLER_0_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08803_ net1093 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[0\] net882 vssd1
+ vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__and3_1
XFILLER_0_147_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09783_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[15\] net788 net783 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06123_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout285_A _07896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11863__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08734_ _05069_ _05070_ _05073_ net703 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__o32a_4
XANTENNA__10620__X _06960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08738__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08665_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[10\] net704 _05001_ _05004_
+ vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__o22ai_4
XANTENNA_fanout452_A _07957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08457__B net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09609__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08596_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[15\] net697 net696 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[15\]
+ _04922_ vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__a221o_1
XANTENNA__14063__B1 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_132_Left_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12694__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout338_X net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08473__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08904__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09217_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[17\] net650 _05532_ _05536_
+ _05538_ vssd1 vssd1 vccd1 vccd1 _05557_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout505_X net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1247_X net1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09148_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[14\] net689 _05459_
+ _05460_ _05475_ vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_72_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09242__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08596__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09079_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] net620 net593 vssd1 vssd1
+ vccd1 vccd1 _05419_ sky130_fd_sc_hd__a21o_1
XANTENNA__12723__A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11110_ _06404_ _06405_ net344 vssd1 vssd1 vccd1 vccd1 _07450_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_9_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_3__f_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_3__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_12090_ net2180 net291 net460 vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_141_Left_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09735__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold770 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2316 sky130_fd_sc_hd__dlygate4sd3_1
X_11041_ _07312_ _07313_ _07380_ vssd1 vssd1 vccd1 vccd1 _07381_ sky130_fd_sc_hd__a21oi_1
Xhold792 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2327 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11773__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14800_ net1282 vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__inv_2
X_15780_ net1197 vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__inv_2
X_12992_ net2841 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[102\] net854 vssd1 vssd1
+ vccd1 vccd1 _02133_ sky130_fd_sc_hd__mux2_1
XANTENNA__08648__A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09848__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1470 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[111\] vssd1 vssd1 vccd1 vccd1
+ net3005 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input13_A DAT_I[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14731_ net1211 vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__inv_2
Xhold1481 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net3016 sky130_fd_sc_hd__dlygate4sd3_1
X_11943_ net2194 net257 net478 vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__mux2_1
Xhold1492 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3027 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09470__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11074__A net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17450_ clknet_leaf_10_wb_clk_i _03137_ _01433_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_14662_ net1228 vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11874_ net1870 net265 net484 vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__mux2_1
X_16401_ clknet_leaf_98_wb_clk_i _02155_ _00384_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[124\]
+ sky130_fd_sc_hd__dfstp_1
X_13613_ team_01_WB.instance_to_wrap.cpu.CU0.bit30 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\]
+ net595 _04053_ vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__a31o_1
X_17381_ clknet_leaf_50_wb_clk_i _03068_ _01364_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10825_ _05618_ net330 vssd1 vssd1 vccd1 vccd1 _07165_ sky130_fd_sc_hd__nor2_1
XFILLER_0_156_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14593_ net1411 vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_45_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16332_ clknet_leaf_120_wb_clk_i _02086_ _00315_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13544_ net986 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] _03995_ _03996_
+ vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_45_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10756_ net335 _07095_ vssd1 vssd1 vccd1 vccd1 _07096_ sky130_fd_sc_hd__nor2_1
XANTENNA__09481__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16263_ clknet_leaf_142_wb_clk_i net1560 _00251_ vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12109__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13475_ _03929_ _03931_ _03935_ vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_97_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10687_ _06888_ _06892_ net533 vssd1 vssd1 vccd1 vccd1 _07027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18002_ net635 vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15214_ net1297 vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12907__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12426_ net3144 net220 net417 vssd1 vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16194_ clknet_leaf_159_wb_clk_i _01954_ _00182_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09233__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10918__A1 _04738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11948__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15145_ net1288 vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__inv_2
XANTENNA__13580__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12357_ _07945_ _07946_ net574 vssd1 vssd1 vccd1 vccd1 _07966_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10394__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09418__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11308_ net721 _07643_ _07646_ vssd1 vssd1 vccd1 vccd1 _07647_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15076_ net1218 vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__inv_2
X_12288_ net2561 net318 net437 vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14027_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[10\] _04253_ _04261_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[114\]
+ _04316_ vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__a221o_1
XANTENNA__11249__A _07588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11239_ _07017_ _07573_ _07578_ _07571_ vssd1 vssd1 vccd1 vccd1 _07579_ sky130_fd_sc_hd__a211oi_4
XANTENNA__09942__A net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_25 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15978_ net1363 vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09839__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14929_ net1423 vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__inv_2
XANTENNA__13183__B net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17717_ clknet_leaf_125_wb_clk_i _03401_ _01658_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10600__B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08450_ net1022 net907 vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__and2_2
X_17648_ clknet_leaf_150_wb_clk_i _03333_ _01589_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14045__B1 _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08381_ _04624_ _04719_ vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__nand2_1
X_17579_ clknet_leaf_96_wb_clk_i _03266_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__dfxtp_1
XANTENNA__12808__A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11712__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08814__A3 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12019__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09002_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[9\] net884 vssd1
+ vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11858__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10909__B2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10499__A_N net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_158_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_158_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08578__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout200_A _07858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10385__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09904_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[5\] net774 _06241_ _06242_
+ _06243_ vssd1 vssd1 vccd1 vccd1 _06244_ sky130_fd_sc_hd__a2111o_1
Xfanout502 _07795_ vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__buf_4
Xfanout513 _05867_ vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09527__B2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout524 net526 vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10137__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17926__1533 vssd1 vssd1 vccd1 vccd1 net1533 _17926__1533/LO sky130_fd_sc_hd__conb_1
XANTENNA_fanout1207_A net1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout535 _05190_ vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__buf_2
XFILLER_0_67_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09852__A net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout546 net547 vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__clkbuf_4
X_09835_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[13\] net749 net745 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06175_ sky130_fd_sc_hd__a22o_1
Xfanout557 net558 vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input5_A DAT_I[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout568 _04520_ vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__buf_2
XANTENNA__12689__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout579 _07752_ vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__buf_2
XANTENNA__10998__A net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout667_A _04801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09766_ _06105_ vssd1 vssd1 vccd1 vccd1 _06106_ sky130_fd_sc_hd__inv_2
XANTENNA__08468__A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08717_ net1097 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[5\] net943 vssd1
+ vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__and3_1
XANTENNA__09290__C net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09697_ net1154 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[21\] net974
+ vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout455_X net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08502__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08648_ net1020 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[10\] net941 vssd1
+ vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__and3_1
XANTENNA__14036__B1 _04266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13821__B net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08579_ _04885_ _04918_ net600 vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__mux2_4
XFILLER_0_3_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10610_ _06948_ _06949_ net540 vssd1 vssd1 vccd1 vccd1 _06950_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08266__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11590_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] _07805_ vssd1 vssd1
+ vccd1 vccd1 _07807_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08634__C net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11341__B _04621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10541_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[31\] net701 _06870_ _06880_
+ vssd1 vssd1 vccd1 vccd1 _06881_ sky130_fd_sc_hd__o22a_2
XFILLER_0_106_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwire947 _04671_ vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__clkbuf_1
XANTENNA__13547__C1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13260_ team_01_WB.instance_to_wrap.cpu.f0.i\[24\] _03751_ vssd1 vssd1 vccd1 vccd1
+ _03752_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_40_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10472_ _06811_ vssd1 vssd1 vccd1 vccd1 _06812_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11768__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12211_ net2653 net226 net443 vssd1 vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13191_ net18 net837 net630 net2026 vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12770__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12142_ net3137 net259 net453 vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__mux2_1
X_12073_ net2318 net267 net460 vssd1 vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__mux2_1
X_16950_ clknet_leaf_12_wb_clk_i _02637_ _00933_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11325__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15901_ net1416 vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__inv_2
X_11024_ _07352_ _07357_ _07363_ vssd1 vssd1 vccd1 vccd1 _07364_ sky130_fd_sc_hd__nand3_1
X_16881_ clknet_leaf_118_wb_clk_i _02568_ _00864_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12599__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12900__B net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15832_ net1339 vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__inv_2
X_15763_ net1198 vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__inv_2
X_12975_ net2850 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[119\] net856 vssd1 vssd1
+ vccd1 vccd1 _02150_ sky130_fd_sc_hd__mux2_1
XANTENNA__12825__B2 _03646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17502_ clknet_leaf_85_wb_clk_i _03189_ _01485_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_14714_ net1191 vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11926_ net3004 net190 net475 vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__mux2_1
X_15694_ net1298 vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__inv_2
XANTENNA__14027__B1 _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17433_ clknet_leaf_71_wb_clk_i _03120_ _01416_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14645_ net1209 vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__inv_2
X_11857_ net1831 net313 net489 vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10808_ _07015_ _07099_ _07146_ _07147_ vssd1 vssd1 vccd1 vccd1 _07148_ sky130_fd_sc_hd__a211o_1
X_17364_ clknet_leaf_22_wb_clk_i _03051_ _01347_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14576_ net1354 vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__inv_2
XANTENNA__09454__B1 _04797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11788_ net2201 net318 net497 vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_136_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13250__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_126_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09002__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16315_ clknet_leaf_119_wb_clk_i _02069_ _00298_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[38\]
+ sky130_fd_sc_hd__dfrtp_1
X_13527_ _03942_ _03981_ vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08662__D1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10739_ _07076_ _07077_ _07078_ vssd1 vssd1 vccd1 vccd1 _07079_ sky130_fd_sc_hd__or3b_1
X_17295_ clknet_leaf_35_wb_clk_i _02982_ _01278_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12915__X _03686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16246_ clknet_leaf_140_wb_clk_i net1734 _00234_ vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_153_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13458_ _03914_ _03915_ _03857_ _03859_ vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__a211o_1
XFILLER_0_152_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11678__S net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12409_ net2492 net254 net420 vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__mux2_1
X_16177_ clknet_leaf_6_wb_clk_i _01937_ _00165_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13389_ _03848_ _03849_ vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__nor2_1
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__buf_2
XANTENNA__12761__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__buf_2
Xoutput127 net127 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput138 net138 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__buf_2
X_15128_ net1213 vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__inv_2
Xoutput149 net149 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
X_15059_ net1394 vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10119__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10314__C net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17662__Q team_01_WB.instance_to_wrap.cpu.DM0.readdata\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17932__1449 vssd1 vssd1 vccd1 vccd1 _17932__1449/HI net1449 sky130_fd_sc_hd__conb_1
XANTENNA__08732__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09620_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[24\] net802 net770 _05958_
+ _05959_ vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12302__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16278__Q team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08719__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09551_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[28\] net757 _05875_ _05879_
+ _05882_ vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12816__A1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12816__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08502_ net1118 net711 net594 vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10827__B1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09482_ net1079 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[30\] net906
+ net688 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[30\] vssd1 vssd1 vccd1
+ vccd1 _05822_ sky130_fd_sc_hd__a32o_1
XFILLER_0_77_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_13__f_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08433_ net1111 _04770_ vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__and2_2
XFILLER_0_93_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08735__B net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout248_A _07842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08364_ _04693_ _04695_ _04700_ _04703_ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__or4_2
XANTENNA__09445__B1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08295_ net1162 net1165 net1167 net1159 vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__nor4b_2
XANTENNA_fanout415_A _03562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13529__C1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1157_A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08751__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13544__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10358__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12752__B1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09285__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08971__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout310 _07931_ vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__clkbuf_2
Xfanout1308 net1309 vssd1 vssd1 vccd1 vccd1 net1308 sky130_fd_sc_hd__buf_4
Xfanout1319 net1321 vssd1 vssd1 vccd1 vccd1 net1319 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout332 _06923_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__clkbuf_2
Xfanout343 _04748_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13816__B net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout354 _03741_ vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__buf_2
XANTENNA_fanout951_A _04662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout365 _03580_ vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__buf_2
Xfanout376 _04969_ vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__clkbuf_4
X_09818_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] _06157_ _04628_ vssd1
+ vssd1 vccd1 vccd1 _06158_ sky130_fd_sc_hd__mux2_4
Xfanout387 _03569_ vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__buf_6
XANTENNA__12212__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout398 _03567_ vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__buf_4
XANTENNA__10521__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_55_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09749_ _06085_ _06086_ _06087_ _06088_ vssd1 vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout837_X net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12760_ net1842 net639 net606 _03601_ vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__a22o_1
XANTENNA__08485__X _04825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08926__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11711_ net718 _07269_ net616 _07905_ vssd1 vssd1 vccd1 vccd1 _07906_ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12691_ net2623 net217 net385 vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14430_ net1335 vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_42_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11642_ net2176 net274 net501 vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13232__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14361_ net1340 vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__inv_2
X_11573_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\] team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\]
+ vssd1 vssd1 vccd1 vccd1 _07790_ sky130_fd_sc_hd__nor2_2
Xinput18 DAT_I[24] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
X_16100_ clknet_leaf_126_wb_clk_i _01875_ _00088_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11794__A1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13312_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[22\] net825 _03791_ _03793_
+ vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__o22a_1
X_17080_ clknet_leaf_49_wb_clk_i _02767_ _01063_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput29 DAT_I[5] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
X_10524_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[31\] net680 _06861_
+ _06862_ _06863_ vssd1 vssd1 vccd1 vccd1 _06864_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_80_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14292_ net1346 vssd1 vssd1 vccd1 vccd1 _00086_ sky130_fd_sc_hd__inv_2
X_16031_ net1325 vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__inv_2
X_13243_ net2988 net354 net350 net1072 vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__a22o_1
XANTENNA__13535__A2 _07600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13279__A team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_150_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10455_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[26\] net822 net805 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06795_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12743__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11546__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13174_ net130 net848 net840 net1938 vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__a22o_1
XANTENNA__09195__C net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10386_ _06723_ _06724_ _06725_ vssd1 vssd1 vccd1 vccd1 _06726_ sky130_fd_sc_hd__or3_1
XFILLER_0_21_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12125_ net2672 net190 net451 vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17982_ net1497 vssd1 vssd1 vccd1 vccd1 la_data_out[24] sky130_fd_sc_hd__buf_2
XANTENNA__13299__A1 _04516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10134__C net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16933_ clknet_leaf_50_wb_clk_i _02620_ _00916_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12056_ net2468 net315 net465 vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__mux2_1
XANTENNA__09923__C net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_9__f_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11007_ _07345_ _07346_ _07344_ vssd1 vssd1 vccd1 vccd1 _07347_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_88_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12122__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16864_ clknet_leaf_46_wb_clk_i _02551_ _00847_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_15815_ net1189 vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__inv_2
X_16795_ clknet_leaf_70_wb_clk_i _02482_ _00778_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14838__A net1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11961__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17910__1521 vssd1 vssd1 vccd1 vccd1 net1521 _17910__1521/LO sky130_fd_sc_hd__conb_1
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15746_ net1315 vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__inv_2
X_12958_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[3\] _05219_ net1039 vssd1
+ vssd1 vccd1 vccd1 _03714_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11909_ net3008 net231 net481 vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15677_ net1311 vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__inv_2
X_12889_ _05704_ net578 net361 vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_28_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14628_ net1387 vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__inv_2
X_17416_ clknet_leaf_62_wb_clk_i _03103_ _01399_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_155_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09427__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17925__1532 vssd1 vssd1 vccd1 vccd1 net1532 _17925__1532/LO sky130_fd_sc_hd__conb_1
X_17347_ clknet_leaf_23_wb_clk_i _03034_ _01330_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12792__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14559_ net1406 vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_151_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09442__A3 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10309__C net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08080_ _04514_ _04528_ _04532_ _04522_ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__o22a_1
XFILLER_0_43_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_wire585_A _05040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17278_ clknet_leaf_84_wb_clk_i _02965_ _01261_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16229_ clknet_leaf_140_wb_clk_i _01989_ _00217_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08290__B net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11537__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08953__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08982_ net1007 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[8\] net911 vssd1
+ vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_149_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_143_Right_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12032__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10512__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09603_ net1145 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[24\] net982
+ vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__and3_1
XFILLER_0_155_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout365_A _03580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11871__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_30_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11724__X _07917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09534_ net996 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[28\] net952 vssd1
+ vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08746__A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09465_ net602 _05803_ _05804_ vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_66_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09418__A0 _05756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08416_ net1116 net1119 net1122 net1125 vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__nor4_2
X_09396_ _05659_ _05681_ _05707_ net560 vssd1 vssd1 vccd1 vccd1 _05736_ sky130_fd_sc_hd__a31o_1
XFILLER_0_148_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10028__A1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08347_ net998 net980 vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12555__X _03566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout418_X net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1062_X net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_102_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_102_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_104_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08278_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[3\] net2086 net1046 vssd1 vssd1
+ vccd1 vccd1 _03409_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13099__A _03719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout999_A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12207__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11528__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10240_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[9\] net747 net737 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06580_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout787_X net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10171_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[10\] net818 net799 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06511_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1105 net1106 vssd1 vssd1 vccd1 vccd1 net1105 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1116 net1117 vssd1 vssd1 vccd1 vccd1 net1116 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1127 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[20\] vssd1 vssd1 vccd1 vccd1
+ net1127 sky130_fd_sc_hd__buf_2
Xfanout1138 net1141 vssd1 vssd1 vccd1 vccd1 net1138 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_35_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout954_X net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1149 net1150 vssd1 vssd1 vccd1 vccd1 net1149 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13150__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11347__A team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13930_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__and2b_2
XANTENNA__10251__A net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout195 _07634_ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11161__C1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10503__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13861_ net1177 net1064 net1660 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[22\]
+ sky130_fd_sc_hd__and3b_1
XANTENNA__11066__B _06158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11781__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15600_ net1272 vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12812_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] net1063 net364 _03636_
+ vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__a22o_1
X_16580_ clknet_leaf_84_wb_clk_i _02267_ _00563_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_69_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13792_ _04165_ _04173_ vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_2_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15531_ net1396 vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__inv_2
X_12743_ net1797 net640 net608 _03589_ vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08375__B _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15462_ net1404 vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12674_ net3126 net286 net390 vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08880__B2 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17201_ clknet_leaf_113_wb_clk_i _02888_ _01184_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_14413_ net1308 vssd1 vssd1 vccd1 vccd1 _00207_ sky130_fd_sc_hd__inv_2
X_11625_ _07836_ _07837_ net612 vssd1 vssd1 vccd1 vccd1 _07838_ sky130_fd_sc_hd__mux2_1
X_15393_ net1278 vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_4_12__f_wb_clk_i_X clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17132_ clknet_leaf_16_wb_clk_i _02819_ _01115_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_14344_ net1330 vssd1 vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__inv_2
X_17931__1448 vssd1 vssd1 vccd1 vccd1 _17931__1448/HI net1448 sky130_fd_sc_hd__conb_1
X_11556_ team_01_WB.instance_to_wrap.cpu.K0.count\[0\] team_01_WB.instance_to_wrap.cpu.K0.enable
+ _07786_ vssd1 vssd1 vccd1 vccd1 _07787_ sky130_fd_sc_hd__and3_1
XFILLER_0_107_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08822__C net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13508__A2 _07056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10507_ _06835_ _06844_ _06845_ _06846_ vssd1 vssd1 vccd1 vccd1 _06847_ sky130_fd_sc_hd__or4_1
X_17063_ clknet_leaf_106_wb_clk_i _02750_ _01046_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12117__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14275_ net1340 vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__inv_2
Xwire585 _05040_ vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__buf_4
X_11487_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[19\] net579 vssd1 vssd1 vccd1
+ vccd1 _07771_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmax_cap329 _05568_ vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16014_ net1329 vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_59_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09188__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13226_ net2808 net352 net348 team_01_WB.instance_to_wrap.cpu.f0.i\[24\] vssd1 vssd1
+ vccd1 vccd1 _01924_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_59_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10438_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[27\] net764 net623 vssd1
+ vssd1 vccd1 vccd1 _06778_ sky130_fd_sc_hd__o21a_1
XANTENNA__11956__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09493__Y _05833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13157_ net1611 net847 _03734_ team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[19\] vssd1
+ vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__a22o_1
X_10369_ _04970_ _05379_ _05494_ _05529_ vssd1 vssd1 vccd1 vccd1 _06709_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_55_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12108_ net2999 net232 net457 vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17965_ net1480 vssd1 vssd1 vccd1 vccd1 la_data_out[7] sky130_fd_sc_hd__buf_2
X_13088_ _03711_ net2987 net853 vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16916_ clknet_leaf_20_wb_clk_i _02603_ _00899_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_12039_ net2498 net236 net463 vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17896_ net1431 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_144_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09950__A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16847_ clknet_leaf_35_wb_clk_i _02534_ _00830_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09648__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16778_ clknet_leaf_32_wb_clk_i _02465_ _00761_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15729_ net1394 vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_0_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_114_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_47_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09250_ _05573_ _05576_ _05587_ _05589_ vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__or4_1
X_08201_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[80\] net3086 net1046 vssd1 vssd1
+ vccd1 vccd1 _03486_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09181_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[16\] net900
+ vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__and3_1
XFILLER_0_145_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10039__C net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11720__A net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08132_ _04488_ team_01_WB.instance_to_wrap.cpu.f0.num\[5\] _04498_ team_01_WB.instance_to_wrap.cpu.f0.i\[2\]
+ _04595_ vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09820__B1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08063_ _04532_ _04539_ vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__nor2_1
XANTENNA__12027__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13856__A_N net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11866__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10194__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1022_A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08965_ net1008 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[8\] net934 vssd1
+ vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout482_A _07949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09563__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08896_ net1107 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[2\] net902 vssd1
+ vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_153_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12697__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1391_A net1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout747_A net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13382__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout368_X net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_8__f_wb_clk_i_X clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_78_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08476__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09103__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08907__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09517_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[29\] net795 _05844_ _05847_
+ _05849_ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13986__A2 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout914_A _04779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09448_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[29\] net681 net659 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[29\]
+ _05787_ vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__a221o_1
XANTENNA__13199__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout702_X net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09379_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[26\] net699 net666 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _05719_ sky130_fd_sc_hd__a22o_1
XANTENNA__12726__A net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08923__B net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11410_ team_01_WB.instance_to_wrap.cpu.f0.i\[20\] _07693_ vssd1 vssd1 vccd1 vccd1
+ _07728_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12390_ _07793_ _07946_ net573 vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__and3_1
XFILLER_0_145_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09811__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09738__C net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08642__C net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11341_ _04511_ _04621_ _07669_ vssd1 vssd1 vccd1 vccd1 _07670_ sky130_fd_sc_hd__and3b_1
X_14060_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[51\] _04236_ _04252_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[107\]
+ vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__a22o_1
X_11272_ _06100_ _06104_ _07089_ vssd1 vssd1 vccd1 vccd1 _07612_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_37_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11776__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13011_ net2336 net1542 net861 vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__mux2_1
X_10223_ _06562_ vssd1 vssd1 vccd1 vccd1 _06563_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_18_Left_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_70_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_30_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input43_A wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09590__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10154_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[11\] net767 _06493_ vssd1
+ vssd1 vccd1 vccd1 _06494_ sky130_fd_sc_hd__o21ba_1
XANTENNA__09473__C net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13123__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14962_ net1266 vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__inv_2
X_17924__1531 vssd1 vssd1 vccd1 vccd1 net1531 _17924__1531/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_7_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17750_ clknet_leaf_118_wb_clk_i _03426_ _01690_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[20\]
+ sky130_fd_sc_hd__dfstp_1
X_10085_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[7\] net797 net730 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06425_ sky130_fd_sc_hd__a22o_1
Xhold7 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[83\] vssd1 vssd1 vccd1 vccd1 net1542
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10412__C net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16701_ clknet_leaf_65_wb_clk_i _02388_ _00684_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13913_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[10\] _04209_ net571 vssd1
+ vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_50_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14893_ net1261 vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__inv_2
X_17681_ clknet_leaf_129_wb_clk_i _03365_ _01622_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_18_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13292__A team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16632_ clknet_leaf_49_wb_clk_i _02319_ _00615_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12400__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13844_ net1179 net1066 net3179 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[5\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_69_241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08817__C net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13775_ team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[1\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\]
+ net605 vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__mux2_1
X_16563_ clknet_leaf_159_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[29\]
+ _00546_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_27_Left_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13977__A2 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10987_ _06313_ _06339_ net551 vssd1 vssd1 vccd1 vccd1 _07327_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_100_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12726_ net1033 team_01_WB.instance_to_wrap.cpu.f0.read_i vssd1 vssd1 vccd1 vccd1
+ _03577_ sky130_fd_sc_hd__nor2_1
X_15514_ net1372 vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__inv_2
X_16494_ clknet_leaf_142_wb_clk_i _02248_ _00477_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15445_ net1277 vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12657_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[29\] net220 net389 vssd1
+ vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11608_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[30\] _07019_ net714 vssd1 vssd1
+ vccd1 vccd1 _07824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08605__A1 net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15376_ net1271 vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__inv_2
XANTENNA__09802__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12588_ _07790_ _07951_ net573 vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__and3_4
XFILLER_0_111_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08552__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17115_ clknet_leaf_71_wb_clk_i _02802_ _01098_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_14327_ net1348 vssd1 vssd1 vccd1 vccd1 _00121_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11539_ net2106 net1174 net590 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] vssd1
+ vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__a22o_1
XANTENNA__10156__A net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14851__A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold407 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1942 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold418 team_01_WB.instance_to_wrap.a1.ADR_I\[31\] vssd1 vssd1 vccd1 vccd1 net1953
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09945__A _06280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17046_ clknet_leaf_28_wb_clk_i _02733_ _01029_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold429 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1964 sky130_fd_sc_hd__dlygate4sd3_1
X_14258_ net1203 vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__inv_2
XANTENNA__14154__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_36_Left_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08908__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13209_ net30 net836 net629 net1601 vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__o22a_1
X_14189_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[14\] _04457_ vssd1 vssd1 vccd1
+ vccd1 _04458_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_74_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout909 _04785_ vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_146_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09581__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15682__A net1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08750_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[4\] net889 vssd1
+ vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__and3_1
Xhold1107 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[105\] vssd1 vssd1 vccd1 vccd1
+ net2642 sky130_fd_sc_hd__dlygate4sd3_1
X_17948_ net1463 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
Xhold1118 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2653 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13665__A1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1129 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 net2664
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08848__X _05188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10322__C net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11676__A0 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09333__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08681_ net1086 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[7\] net882 vssd1
+ vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__and3_1
X_17879_ clknet_leaf_135_wb_clk_i _03554_ _01819_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12310__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08296__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_max_cap967_X net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09302_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[22\] net904
+ vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__and3_1
XFILLER_0_152_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09233_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[21\] net686 net682 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[21\]
+ _05571_ vssd1 vssd1 vccd1 vccd1 _05573_ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10618__X _06958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout230_A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09164_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[16\] net904
+ vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__and3_1
XFILLER_0_146_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08115_ team_01_WB.instance_to_wrap.cpu.f0.i\[1\] team_01_WB.instance_to_wrap.cpu.f0.num\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08462__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13929__X _04221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15857__A net1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09095_ net1093 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[13\] net892
+ vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1237_A net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08046_ net1633 net569 _04526_ team_01_WB.instance_to_wrap.cpu.f0.i\[9\] vssd1 vssd1
+ vccd1 vccd1 _03545_ sky130_fd_sc_hd__a22o_1
Xclkbuf_4_2__f_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_2__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__14145__A2 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold930 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[42\] vssd1 vssd1 vccd1 vccd1
+ net2465 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold941 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2476 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout697_A net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09557__C1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold952 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold963 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold974 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2509 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10167__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1404_A net1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold985 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2520 sky130_fd_sc_hd__dlygate4sd3_1
Xhold996 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2531 sky130_fd_sc_hd__dlygate4sd3_1
X_09997_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[2\] _04678_ _06333_
+ _06334_ _06336_ vssd1 vssd1 vccd1 vccd1 _06337_ sky130_fd_sc_hd__a2111o_2
XANTENNA__09293__C net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout864_A net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout485_X net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15592__A net1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08948_ net1027 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[6\] net890 vssd1
+ vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_4_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1630 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net3165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1641 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1 net3176
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09324__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13824__B net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08879_ _05211_ _05215_ _05218_ net704 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__o32a_4
Xhold1652 team_01_WB.instance_to_wrap.cpu.c0.count\[13\] vssd1 vssd1 vccd1 vccd1 net3187
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout652_X net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17930__1447 vssd1 vssd1 vccd1 vccd1 _17930__1447/HI net1447 sky130_fd_sc_hd__conb_1
XANTENNA__11184__X _07524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10910_ _07054_ _07235_ _07241_ _07249_ vssd1 vssd1 vccd1 vccd1 _07250_ sky130_fd_sc_hd__a31o_1
XANTENNA__12220__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11890_ net2062 net315 net485 vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__mux2_1
XANTENNA__08637__C net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10841_ _06065_ _06098_ _06636_ _06671_ net549 net538 vssd1 vssd1 vccd1 vccd1 _07181_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11344__B team_01_WB.instance_to_wrap.cpu.f0.i\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_39_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout917_X net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13560_ net720 _07171_ net1073 vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__o21a_1
XFILLER_0_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10772_ _06598_ _06604_ _06742_ vssd1 vssd1 vccd1 vccd1 _07112_ sky130_fd_sc_hd__a21o_1
X_12511_ net1994 net249 net410 vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__mux2_1
XANTENNA__10642__A1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13491_ _03841_ _03842_ _03950_ _03839_ vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__a31o_1
XFILLER_0_109_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15230_ net1345 vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12442_ net2188 net256 net416 vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15161_ net1235 vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__inv_2
X_12373_ net1894 net261 net424 vssd1 vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12890__S net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10945__A2 _06188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14112_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[38\] _04230_ _04259_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09765__A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11324_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[2\] team_01_WB.instance_to_wrap.cpu.DM0.data_i\[1\]
+ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[0\] _07658_ vssd1 vssd1 vccd1 vccd1
+ _07659_ sky130_fd_sc_hd__or4_1
XANTENNA__14136__A2 _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15092_ net1399 vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_95_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14043_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[3\] _04249_ _04255_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[115\]
+ _04331_ vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__a221o_1
X_11255_ net523 _07534_ _07594_ vssd1 vssd1 vccd1 vccd1 _07595_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10158__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10206_ net1143 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[8\] net955 vssd1
+ vssd1 vccd1 vccd1 _06546_ sky130_fd_sc_hd__and3_1
XANTENNA__11519__B net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11186_ _07234_ _07483_ net525 vssd1 vssd1 vccd1 vccd1 _07526_ sky130_fd_sc_hd__mux2_1
X_17802_ clknet_leaf_122_wb_clk_i net2946 _01742_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[72\]
+ sky130_fd_sc_hd__dfrtp_1
X_10137_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[11\] net807 net782 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06477_ sky130_fd_sc_hd__a22o_1
XANTENNA__13647__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15994_ net1353 vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__inv_2
XANTENNA__09315__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11658__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17733_ clknet_leaf_125_wb_clk_i _03409_ _01673_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10068_ _06285_ _06407_ vssd1 vssd1 vccd1 vccd1 _06408_ sky130_fd_sc_hd__nand2_1
X_14945_ net1280 vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_141_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12130__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17664_ clknet_leaf_0_wb_clk_i _03349_ _01605_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14876_ net1243 vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__inv_2
XANTENNA__09005__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_56 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10881__A1 _05566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08547__C net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16615_ clknet_leaf_105_wb_clk_i _02302_ _00598_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13827_ net2608 net831 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[20\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__09079__A1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17595_ clknet_leaf_89_wb_clk_i _03282_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13758_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[13\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[12\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[14\] vssd1 vssd1 vccd1 vccd1 _04147_
+ sky130_fd_sc_hd__or3b_1
X_16546_ clknet_leaf_2_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[12\]
+ _00529_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12709_ net2172 net249 net386 vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13689_ team_01_WB.instance_to_wrap.cpu.c0.count\[6\] team_01_WB.instance_to_wrap.cpu.c0.count\[5\]
+ team_01_WB.instance_to_wrap.cpu.c0.count\[15\] team_01_WB.instance_to_wrap.cpu.c0.count\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__or4bb_1
X_16477_ clknet_leaf_141_wb_clk_i _02231_ _00460_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15428_ net1222 vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11189__A2 _07527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_44_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15359_ net1312 vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold204 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1739 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09675__A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold215 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1750 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14127__A2 _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold226 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net1761 sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1772 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09920_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[4\] net808 net772 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06260_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_113_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold248 _03529_ vssd1 vssd1 vccd1 vccd1 net1783 sky130_fd_sc_hd__dlygate4sd3_1
X_17029_ clknet_leaf_46_wb_clk_i _02716_ _01012_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold259 net131 vssd1 vssd1 vccd1 vccd1 net1794 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12305__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10149__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout706 net708 vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout717 _04723_ vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__buf_2
X_09851_ _05454_ _06190_ vssd1 vssd1 vccd1 vccd1 _06191_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09554__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout728 _04720_ vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__clkbuf_4
Xfanout739 net741 vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__buf_6
X_08802_ net1011 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[0\] net879 vssd1
+ vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__and3_1
X_09782_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[15\] net820 _06120_
+ _06121_ vssd1 vssd1 vccd1 vccd1 _06122_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13638__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08578__X _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08733_ _05061_ _05064_ _05071_ _05072_ vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__or4_1
XANTENNA__09306__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_53_Left_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08664_ _04995_ _04996_ _05002_ _05003_ vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__or4_1
XANTENNA__12040__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08595_ _04932_ _04933_ _04934_ vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout445_A _07959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10624__A1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout612_A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08473__B net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1354_A net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09216_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[17\] net654 _05535_
+ _05542_ _05553_ vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09288__C net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17923__1530 vssd1 vssd1 vccd1 vccd1 net1530 _17923__1530/LO sky130_fd_sc_hd__conb_1
X_09147_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[14\] net681 _05467_
+ _05472_ net707 vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_20_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15587__A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout400_X net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12916__A3 _03686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08045__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09242__A1 net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10388__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10927__A2 _07227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14118__A2 _04246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13819__B net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09078_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] net620 _04845_ vssd1 vssd1
+ vccd1 vccd1 _05418_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout981_A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12723__B team_01_WB.instance_to_wrap.cpu.f0.write_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08029_ team_01_WB.instance_to_wrap.cpu.f0.state\[7\] net569 vssd1 vssd1 vccd1 vccd1
+ _04525_ sky130_fd_sc_hd__nor2_2
XANTENNA__12215__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold760 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2306 sky130_fd_sc_hd__dlygate4sd3_1
Xhold782 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2317 sky130_fd_sc_hd__dlygate4sd3_1
X_11040_ _07295_ _07296_ vssd1 vssd1 vccd1 vccd1 _07380_ sky130_fd_sc_hd__nor2_1
XANTENNA__09545__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold793 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[9\] vssd1 vssd1 vccd1 vccd1 net2328
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout867_X net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13629__A1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12991_ net2477 net2337 net858 vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__mux2_1
Xhold1460 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2995 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08505__B1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11104__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1471 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 net3006
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14730_ net1210 vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__inv_2
X_11942_ net2648 net232 net477 vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__mux2_1
Xhold1482 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net3017 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10312__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1493 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net3028 sky130_fd_sc_hd__dlygate4sd3_1
X_14661_ net1305 vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__inv_2
XANTENNA__10863__B2 _06920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11873_ net1814 net233 net483 vssd1 vssd1 vccd1 vccd1 _03105_ sky130_fd_sc_hd__mux2_1
X_13612_ _03888_ _04052_ vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__and2b_1
XFILLER_0_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16400_ clknet_leaf_95_wb_clk_i net1789 _00383_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[123\]
+ sky130_fd_sc_hd__dfrtp_1
X_10824_ _05619_ net507 vssd1 vssd1 vccd1 vccd1 _07164_ sky130_fd_sc_hd__nand2_1
X_17380_ clknet_leaf_84_wb_clk_i _03067_ _01363_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14592_ net1353 vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13543_ net720 _07111_ net1073 vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__o21a_1
X_16331_ clknet_leaf_117_wb_clk_i _02085_ _00314_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[54\]
+ sky130_fd_sc_hd__dfrtp_1
X_10755_ _04844_ net510 vssd1 vssd1 vccd1 vccd1 _07095_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_45_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08383__B team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_923 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10091__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16262_ clknet_leaf_152_wb_clk_i net1586 _00250_ vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__dfrtp_1
X_13474_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] _05592_ _05616_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_97_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09198__C net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10686_ _06979_ _07025_ vssd1 vssd1 vccd1 vccd1 _07026_ sky130_fd_sc_hd__nand2_1
X_18001_ net636 vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__clkbuf_1
X_15213_ net1268 vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__inv_2
XANTENNA__13565__B1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12425_ net2520 net221 net415 vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16193_ clknet_leaf_159_wb_clk_i _01953_ _00181_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10379__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15144_ net1376 vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__inv_2
X_12356_ net2220 net289 net428 vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09784__A2 _04634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11307_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] _05116_ vssd1 vssd1 vccd1
+ vccd1 _07646_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08830__C net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15075_ net1220 vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__inv_2
X_12287_ net1971 net306 net438 vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__mux2_1
XANTENNA__12125__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14026_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[98\] _04244_ _04258_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[58\]
+ vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__a22o_1
X_11238_ net553 _07266_ _07572_ _07575_ _07577_ vssd1 vssd1 vccd1 vccd1 _07578_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09536__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11964__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10777__S1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10551__A0 _06707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11169_ _07269_ _07290_ _07308_ _07508_ vssd1 vssd1 vccd1 vccd1 _07509_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_101_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10570__A_N _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15977_ net1403 vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17716_ clknet_leaf_125_wb_clk_i _03400_ _01657_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_14928_ net1274 vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_69_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10303__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12795__S net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17647_ clknet_leaf_150_wb_clk_i _03332_ _01588_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14859_ net1397 vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08380_ _04624_ _04719_ vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17578_ clknet_leaf_95_wb_clk_i _03265_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17669__CLK clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16529_ clknet_leaf_0_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[27\]
+ _00512_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10082__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09001_ net1095 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[9\] net904 vssd1
+ vssd1 vccd1 vccd1 _05341_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_115_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09224__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[17\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15200__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09775__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08740__C net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13308__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12035__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09692__X _06032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09903_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[5\] net816 net743 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06243_ sky130_fd_sc_hd__a22o_1
Xfanout503 _06857_ vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__buf_4
Xfanout514 net515 vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__clkbuf_4
Xfanout525 net526 vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11874__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout536 net538 vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout395_A _03567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09834_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[13\] net801 net769 vssd1
+ vssd1 vccd1 vccd1 _06174_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_127_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_127_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout547 _05152_ vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__buf_2
XANTENNA__10542__A0 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1102_A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout558 _05114_ vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08749__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10998__B _05263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout569 net570 vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__clkbuf_4
X_09765_ net507 _06099_ vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09571__C net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout562_A net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08468__B net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08716_ net1017 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[5\] net932 vssd1
+ vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__and3_1
X_09696_ _06034_ _06035_ vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__or2_1
X_08647_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[10\] net889
+ vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout448_X net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout827_A _04579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13390__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08578_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[19\] net701 _04900_ _04917_
+ vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__o22a_4
XFILLER_0_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09463__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout615_X net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10540_ _06875_ _06877_ _06878_ _06879_ vssd1 vssd1 vccd1 vccd1 _06880_ sky130_fd_sc_hd__or4_1
XFILLER_0_146_271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10471_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] net627 _06809_ _06810_
+ vssd1 vssd1 vccd1 vccd1 _06811_ sky130_fd_sc_hd__a22o_4
XFILLER_0_17_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12210_ net2564 net285 net446 vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13190_ net19 net835 net628 net1643 vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__o22a_1
XFILLER_0_121_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout984_X net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08650__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12770__A1 _07135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12141_ net3114 net231 net453 vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__mux2_1
XANTENNA__10254__A net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09518__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12072_ net1941 net234 net459 vssd1 vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__mux2_1
Xhold590 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2125 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11784__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11023_ _07361_ _07362_ _07223_ _07359_ vssd1 vssd1 vccd1 vccd1 _07363_ sky130_fd_sc_hd__a211oi_1
X_15900_ net1360 vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10541__X _06881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16880_ clknet_leaf_109_wb_clk_i _02567_ _00863_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10533__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15831_ net1339 vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__inv_2
XANTENNA__08378__B _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15762_ net1198 vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__inv_2
X_12974_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[112\] net1981 net852 vssd1 vssd1
+ vccd1 vccd1 _02151_ sky130_fd_sc_hd__mux2_1
XANTENNA__09151__A0 _05456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16566__CLK clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10420__C net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1290 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2825 sky130_fd_sc_hd__dlygate4sd3_1
X_17501_ clknet_leaf_65_wb_clk_i _03188_ _01484_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_14713_ net1188 vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11925_ _07790_ net575 _07946_ vssd1 vssd1 vccd1 vccd1 _07950_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_86_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15693_ net1263 vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08665__Y _05005_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17432_ clknet_leaf_49_wb_clk_i _03119_ _01415_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11856_ net2300 net317 net490 vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__mux2_1
X_14644_ net1244 vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10807_ _07004_ _07100_ net327 _06988_ vssd1 vssd1 vccd1 vccd1 _07147_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_64_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08825__C net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17363_ clknet_leaf_18_wb_clk_i _03050_ _01346_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_14575_ net1406 vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_136_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11787_ net1779 net306 net497 vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16314_ clknet_leaf_100_wb_clk_i _02068_ _00297_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[37\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10738_ _06964_ _07055_ _07068_ net528 vssd1 vssd1 vccd1 vccd1 _07078_ sky130_fd_sc_hd__a211o_1
X_13526_ _03851_ _03852_ vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17294_ clknet_leaf_36_wb_clk_i _02981_ _01277_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_79 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13457_ _03859_ _03917_ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__or2_1
X_16245_ clknet_leaf_142_wb_clk_i net1623 _00233_ vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_153_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10669_ _07006_ _07008_ net541 vssd1 vssd1 vccd1 vccd1 _07009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12408_ net2984 net259 net421 vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__mux2_1
XANTENNA__09757__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13388_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] _05727_ vssd1 vssd1
+ vccd1 vccd1 _03849_ sky130_fd_sc_hd__nor2_1
X_16176_ clknet_leaf_6_wb_clk_i _01936_ _00164_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__buf_2
XANTENNA__12761__A1 _07154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__buf_2
X_12339_ net2985 net266 net427 vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_110_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput128 net128 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__buf_2
X_15127_ net1243 vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__inv_2
XANTENNA__10164__A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput139 net139 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__buf_2
XFILLER_0_142_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15058_ net1290 vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__inv_2
XANTENNA__11694__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14009_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[121\] _04250_ _04297_ _04299_
+ vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__a211o_1
XANTENNA__09390__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_108_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_20_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09550_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[28\] net795 _05873_ _05877_
+ _05878_ vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_108_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08501_ _04717_ _04752_ _04838_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1
+ vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__o31a_2
XANTENNA__10827__A1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09481_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[30\] net698 net696 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _05821_ sky130_fd_sc_hd__a22o_1
XANTENNA__12819__A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08432_ net1026 net931 vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__and2_2
XFILLER_0_65_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08735__C net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08363_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[30\] net738 _04701_
+ _04702_ net768 vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_19_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09445__A1 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10339__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09996__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08294_ net1154 net979 vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__and2_4
XFILLER_0_116_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11869__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout310_A _07931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout408_A _03564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1052_A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09748__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09566__C net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12752__A1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12752__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1317_A net1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout300 net303 vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__buf_2
Xfanout311 _07931_ vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__buf_2
XANTENNA_fanout777_A _04666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout398_X net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1309 net1310 vssd1 vssd1 vccd1 vccd1 net1309 sky130_fd_sc_hd__buf_2
XFILLER_0_100_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout333 net334 vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10802__A _05657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout344 _04748_ vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__clkbuf_2
Xfanout355 _03741_ vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout366 _07759_ vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09381__B1 _04797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09920__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09817_ _06149_ _06153_ _06155_ _06156_ vssd1 vssd1 vccd1 vccd1 _06157_ sky130_fd_sc_hd__o31a_2
Xfanout377 _04750_ vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__clkbuf_4
Xfanout388 _03569_ vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__clkbuf_4
Xfanout399 _03566_ vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__buf_8
XFILLER_0_154_1012 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09748_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[20\] net802 _06070_
+ _06078_ _06080_ vssd1 vssd1 vccd1 vccd1 _06088_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_115_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13832__B net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout732_X net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09679_ _06016_ _06017_ _06018_ vssd1 vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__or3_1
XANTENNA__08487__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11710_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[9\] net714 vssd1 vssd1 vccd1
+ vccd1 _07905_ sky130_fd_sc_hd__or2_1
XANTENNA__08926__B net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_95_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12690_ net2421 net219 net385 vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08645__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_24_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11641_ _07848_ _07849_ _07850_ net611 vssd1 vssd1 vccd1 vccd1 _07851_ sky130_fd_sc_hd__a22o_2
XFILLER_0_154_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14944__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10046__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14360_ net1336 vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__inv_2
XANTENNA__09987__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11572_ _04726_ _04752_ net620 vssd1 vssd1 vccd1 vccd1 _07789_ sky130_fd_sc_hd__or3_1
XANTENNA__08942__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13311_ net564 _07709_ _03792_ net828 vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__a31o_1
XANTENNA__11779__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput19 DAT_I[25] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
X_10523_ net1003 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[31\] net929 vssd1
+ vssd1 vccd1 vccd1 _06863_ sky130_fd_sc_hd__and3_1
X_14291_ net1346 vssd1 vssd1 vccd1 vccd1 _00085_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16030_ net1323 vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__inv_2
X_13242_ net2485 net355 net351 team_01_WB.instance_to_wrap.cpu.f0.i\[8\] vssd1 vssd1
+ vccd1 vccd1 _01908_ sky130_fd_sc_hd__a22o_1
XANTENNA_input73_A wbs_stb_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10454_ net1148 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[26\] net982
+ vssd1 vssd1 vccd1 vccd1 _06794_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13173_ net133 net848 net840 net1874 vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__a22o_1
X_10385_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[16\] net759 net736 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06725_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12751__X _03595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12124_ _07791_ net575 _07793_ vssd1 vssd1 vccd1 vccd1 _07957_ sky130_fd_sc_hd__and3_4
XANTENNA__10415__C net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17981_ net1496 vssd1 vssd1 vccd1 vccd1 la_data_out[23] sky130_fd_sc_hd__buf_2
XFILLER_0_20_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11367__X _07696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12055_ net1965 net319 net466 vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__mux2_1
X_16932_ clknet_leaf_84_wb_clk_i _02619_ _00915_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12403__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10506__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11006_ _05729_ _06812_ vssd1 vssd1 vccd1 vccd1 _07346_ sky130_fd_sc_hd__nor2_1
XANTENNA__09372__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16863_ clknet_leaf_45_wb_clk_i _02550_ _00846_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_15814_ net1205 vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__inv_2
X_16794_ clknet_leaf_76_wb_clk_i _02481_ _00777_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13742__B net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15745_ net1280 vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__inv_2
X_12957_ net1656 net870 net357 _03713_ vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_104_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11908_ net2080 net261 net480 vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10285__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15676_ net1245 vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__inv_2
X_12888_ net1609 net869 net356 _03666_ vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__a22o_1
XANTENNA__09013__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17415_ clknet_leaf_107_wb_clk_i _03102_ _01398_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_155_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14627_ net1381 vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11839_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[19\] net238 net487 vssd1
+ vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_155_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11234__A1 _04738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17346_ clknet_leaf_56_wb_clk_i _03033_ _01329_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09948__A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14558_ net1401 vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11689__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13509_ _03966_ _03967_ net1074 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__o2bb2a_1
X_17277_ clknet_leaf_64_wb_clk_i _02964_ _01260_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_14489_ net1364 vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14184__B1 net1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16228_ clknet_leaf_140_wb_clk_i net1619 _00216_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10606__B _06250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13757__X _04146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12734__B2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16159_ clknet_leaf_134_wb_clk_i _01922_ _00147_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10745__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08998__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10325__C net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08981_ net1088 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[8\] net904 vssd1
+ vssd1 vccd1 vccd1 _05321_ sky130_fd_sc_hd__and3_1
XANTENNA__17673__Q team_01_WB.instance_to_wrap.cpu.DM0.readdata\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12313__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09902__A2 _04654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_143_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_138_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_127_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09602_ net1146 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[24\] net979
+ vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09533_ net1152 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[28\] net982
+ vssd1 vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout260_A _07888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout358_A net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09464_ net598 _05802_ vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__or2_1
XANTENNA__10276__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08415_ net711 _04751_ _04752_ vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08465__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09395_ _05659_ _05681_ net560 vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08346_ net1143 net945 vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08277_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[4\] net1538 net1042 vssd1 vssd1
+ vccd1 vccd1 _03410_ sky130_fd_sc_hd__mux2_1
XANTENNA__10984__A0 _07277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08481__B net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09296__C net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout894_A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11528__A2 net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15595__A net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_142_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_142_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_132_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10170_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[10\] net806 net771 vssd1
+ vssd1 vccd1 vccd1 _06510_ sky130_fd_sc_hd__a21o_1
XANTENNA__13827__B net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout682_X net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11187__X _07527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11628__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1106 net1114 vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__clkbuf_2
Xfanout1117 net1118 vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1128 net1129 vssd1 vssd1 vccd1 vccd1 net1128 sky130_fd_sc_hd__clkbuf_2
Xfanout1139 net1141 vssd1 vssd1 vccd1 vccd1 net1139 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_35_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09354__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08002__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout185 net186 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_4
Xfanout196 _07633_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__clkbuf_4
X_13860_ net1181 net1065 net3178 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[21\]
+ sky130_fd_sc_hd__and3b_1
X_12811_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[6\] _07323_ net1037 vssd1 vssd1
+ vccd1 vccd1 _03636_ sky130_fd_sc_hd__mux2_1
XANTENNA__13989__B1 _04254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13791_ _01834_ _01833_ vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_2_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11363__A team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15530_ net1385 vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__inv_2
X_12742_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] net1062 net364 _03588_
+ vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12673_ net2657 net254 net388 vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__mux2_1
X_15461_ net1286 vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13205__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11650__X _07858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17200_ clknet_leaf_21_wb_clk_i _02887_ _01183_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10019__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11624_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] _07819_ vssd1 vssd1
+ vccd1 vccd1 _07837_ sky130_fd_sc_hd__xor2_1
X_14412_ net1359 vssd1 vssd1 vccd1 vccd1 _00206_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15392_ net1272 vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12964__A1 _05150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17131_ clknet_leaf_11_wb_clk_i _02818_ _01114_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_14343_ net1338 vssd1 vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__inv_2
X_11555_ net1182 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.next_state
+ sky130_fd_sc_hd__inv_2
XFILLER_0_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10506_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[31\] net815 net806 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06846_ sky130_fd_sc_hd__a22o_1
X_17062_ clknet_leaf_72_wb_clk_i _02749_ _01045_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14274_ net1340 vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11486_ net367 _07770_ net1924 net875 vssd1 vssd1 vccd1 vccd1 _03351_ sky130_fd_sc_hd__o2bb2a_1
X_13225_ net2936 net353 net349 team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1
+ vccd1 vccd1 _01925_ sky130_fd_sc_hd__a22o_1
X_16013_ net1348 vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_59_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10437_ _06766_ _06768_ _06773_ _06776_ vssd1 vssd1 vccd1 vccd1 _06777_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_59_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13156_ net120 net846 net839 net1641 vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__a22o_1
X_10368_ _06707_ vssd1 vssd1 vccd1 vccd1 _06708_ sky130_fd_sc_hd__inv_2
X_12107_ net2221 net264 net456 vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__mux2_1
X_17964_ net1479 vssd1 vssd1 vccd1 vccd1 la_data_out[6] sky130_fd_sc_hd__buf_2
XANTENNA__10442__A net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13087_ _03710_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[7\] net852 vssd1 vssd1
+ vccd1 vccd1 _02038_ sky130_fd_sc_hd__mux2_1
XANTENNA__12133__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10299_ net505 _06638_ vssd1 vssd1 vccd1 vccd1 _06639_ sky130_fd_sc_hd__nand2_1
XANTENNA__09008__A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12038_ net2107 net239 net463 vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__mux2_1
X_16915_ clknet_leaf_18_wb_clk_i _02602_ _00898_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_17895_ net1517 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
XFILLER_0_109_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11972__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16846_ clknet_leaf_28_wb_clk_i _02533_ _00829_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_144_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16134__CLK clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17969__1484 vssd1 vssd1 vccd1 vccd1 _17969__1484/HI net1484 sky130_fd_sc_hd__conb_1
XFILLER_0_88_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16777_ clknet_leaf_40_wb_clk_i _02464_ _00760_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13989_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[72\] _04235_ _04254_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[96\]
+ _04271_ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_122_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15728_ net1275 vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15659_ net1398 vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__inv_2
XANTENNA__08871__A2 _04800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08200_ net2799 net2864 net1057 vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__mux2_1
X_09180_ net1091 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[16\] net892
+ vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__and3_1
XANTENNA__11207__B2 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13601__C1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08582__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16572__Q team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08131_ _04465_ team_01_WB.instance_to_wrap.cpu.f0.num\[31\] team_01_WB.instance_to_wrap.cpu.f0.num\[26\]
+ _04469_ _04588_ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__a221o_1
XANTENNA__11720__B _07308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17329_ clknet_leaf_117_wb_clk_i _03016_ _01312_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12308__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09820__A1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08623__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08062_ _04513_ team_01_WB.instance_to_wrap.cpu.K0.code\[1\] team_01_WB.instance_to_wrap.cpu.K0.code\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__or3b_2
XANTENNA__10430__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_1__f_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_1__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13928__A team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12043__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08964_ net1087 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[8\] net896 vssd1
+ vssd1 vccd1 vccd1 _05304_ sky130_fd_sc_hd__and3_1
XANTENNA__08139__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09336__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13934__Y _04226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08895_ net1025 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[2\] net907 vssd1
+ vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__and3_1
XANTENNA__11882__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout475_A _07950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11735__X _07926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10497__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08757__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12891__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13382__B _05803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout642_A net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1384_A net1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10249__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11446__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09516_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[29\] net812 net770 _05840_
+ _05843_ vssd1 vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_116_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09447_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[29\] net673 net647 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout430_X net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1172_X net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout907_A net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09378_ _05716_ _05717_ vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12726__B team_01_WB.instance_to_wrap.cpu.f0.read_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12946__A1 _05337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08329_ net993 net957 vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__and2_1
XANTENNA__12218__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10957__A0 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09272__C1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08614__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09875__X _06215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11340_ _07651_ team_01_WB.instance_to_wrap.cpu.f0.state\[6\] _04576_ vssd1 vssd1
+ vccd1 vccd1 _07669_ sky130_fd_sc_hd__or3b_1
XANTENNA__14148__B1 _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout897_X net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11271_ _07601_ _07602_ _07610_ vssd1 vssd1 vccd1 vccd1 _07611_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_37_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13010_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[76\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[84\]
+ net855 vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10222_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] net625 _06560_ _06561_
+ vssd1 vssd1 vccd1 vccd1 _06562_ sky130_fd_sc_hd__a22o_4
XANTENNA__09575__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10153_ _06486_ _06490_ _06492_ vssd1 vssd1 vccd1 vccd1 _06493_ sky130_fd_sc_hd__nor3_1
XANTENNA__09327__B1 _04808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11077__B _04919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10084_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[7\] net793 net748 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06424_ sky130_fd_sc_hd__a22o_1
X_14961_ net1394 vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_7_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input36_A gpio_in[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14669__A net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11792__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 _02122_ vssd1 vssd1 vccd1 vccd1 net1543 sky130_fd_sc_hd__dlygate4sd3_1
X_16700_ clknet_leaf_58_wb_clk_i _02387_ _00683_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13912_ _04209_ net571 _04208_ vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_50_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17680_ clknet_leaf_129_wb_clk_i _03364_ _01621_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_14892_ net1260 vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__inv_2
XANTENNA__12882__B1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16631_ clknet_leaf_14_wb_clk_i _02318_ _00614_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13843_ net1180 net1067 net3174 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[4\]
+ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_18_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11093__A net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11437__A1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16562_ clknet_leaf_157_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[28\]
+ _00545_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13774_ team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[0\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[0\]
+ _04146_ vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__mux2_1
X_10986_ _07012_ _07325_ net541 vssd1 vssd1 vccd1 vccd1 _07326_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15513_ net1239 vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__inv_2
X_12725_ team_01_WB.instance_to_wrap.cpu.DM0.state\[0\] _07783_ team_01_WB.instance_to_wrap.cpu.DM0.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_139_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16493_ clknet_leaf_152_wb_clk_i _02247_ _00476_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12917__A _05564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09498__A _04706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15444_ net1399 vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12656_ net2848 net222 net387 vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08833__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11607_ net2530 net191 net499 vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__mux2_1
X_15375_ net1391 vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__inv_2
X_12587_ net1947 net290 net400 vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__mux2_1
XANTENNA__12128__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17114_ clknet_leaf_79_wb_clk_i _02801_ _01097_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14139__B1 _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14326_ net1331 vssd1 vssd1 vccd1 vccd1 _00120_ sky130_fd_sc_hd__inv_2
X_11538_ net2146 net1174 net590 net1168 vssd1 vssd1 vccd1 vccd1 _03314_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold408 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1943 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11967__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold419 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1954 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17045_ clknet_leaf_112_wb_clk_i _02732_ _01028_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_14257_ net1206 vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__inv_2
X_11469_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[28\] net579 vssd1 vssd1 vccd1
+ vccd1 _07762_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13208_ net31 net836 net629 net2158 vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__o22a_1
X_14188_ net1427 _04456_ _04457_ vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_74_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09664__C net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_146_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13139_ net101 net844 net633 net1569 vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_146_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17947_ net1462 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
Xhold1108 _02144_ vssd1 vssd1 vccd1 vccd1 net2643 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12798__S net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1119 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2654 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14579__A net1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13665__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08680_ net1006 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[7\] net926 vssd1
+ vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__and3_1
XANTENNA__11676__A1 _07541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12873__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17878_ clknet_leaf_135_wb_clk_i _03553_ _01818_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16567__Q team_01_WB.instance_to_wrap.cpu.DM0.ihit vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08541__B2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16829_ clknet_leaf_65_wb_clk_i _02516_ _00812_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08296__B net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09301_ net1005 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[22\] net904
+ vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14090__A2 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08844__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09232_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[21\] net691 net685 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08743__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09201__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12928__A1 _05490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09163_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[16\] net654 _05500_
+ _05501_ _05502_ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_8_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12038__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10347__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08114_ team_01_WB.instance_to_wrap.cpu.f0.i\[11\] team_01_WB.instance_to_wrap.cpu.f0.num\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__xnor2_1
X_09094_ net1011 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[13\] net918 vssd1
+ vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__and3_1
XANTENNA__11877__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08045_ net1565 net570 net346 team_01_WB.instance_to_wrap.cpu.f0.i\[10\] vssd1 vssd1
+ vccd1 vccd1 _03546_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold920 _03524_ vssd1 vssd1 vccd1 vccd1 net2455 sky130_fd_sc_hd__dlygate4sd3_1
Xhold931 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2466 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1132_A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold942 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[95\] vssd1 vssd1 vccd1 vccd1
+ net2477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold953 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2488 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold964 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2499 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09574__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold975 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2510 sky130_fd_sc_hd__dlygate4sd3_1
Xhold986 team_01_WB.instance_to_wrap.cpu.f0.num\[2\] vssd1 vssd1 vccd1 vccd1 net2521
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08765__D1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15873__A net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold997 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[107\] vssd1 vssd1 vccd1 vccd1
+ net2532 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13096__C net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09996_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[2\] net762 _06317_ _06335_
+ vssd1 vssd1 vccd1 vccd1 _06336_ sky130_fd_sc_hd__a211o_1
X_08947_ net1111 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[6\] net943 vssd1
+ vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout380_X net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout478_X net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout857_A net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1620 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[28\] vssd1 vssd1 vccd1 vccd1
+ net3155 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11667__A1 _07251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1631 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net3166 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10810__A net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1642 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 net3177
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12501__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08878_ _05208_ _05212_ _05216_ _05217_ vssd1 vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__or4_1
Xhold1653 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 net3188
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1387_X net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10840_ net374 _06158_ _06707_ net371 net550 net535 vssd1 vssd1 vccd1 vccd1 _07180_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_79_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14081__A2 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10771_ net562 _07092_ _07093_ _07110_ vssd1 vssd1 vccd1 vccd1 _07111_ sky130_fd_sc_hd__a31o_2
XANTENNA_fanout812_X net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08835__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12510_ net2791 net227 net407 vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__mux2_1
X_13490_ _03842_ _03950_ vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08653__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12441_ net2038 net258 net418 vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09796__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13592__A1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12372_ net2748 net265 net424 vssd1 vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__mux2_1
X_15160_ net1212 vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__inv_2
XANTENNA__09260__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11787__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10945__A3 _06216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11323_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[7\] team_01_WB.instance_to_wrap.cpu.DM0.data_i\[6\]
+ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[5\] team_01_WB.instance_to_wrap.cpu.DM0.data_i\[3\]
+ vssd1 vssd1 vccd1 vccd1 _07658_ sky130_fd_sc_hd__or4_1
X_14111_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[102\] _04244_ _04247_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[70\]
+ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__a22o_1
X_15091_ net1405 vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__inv_2
X_17968__1483 vssd1 vssd1 vccd1 vccd1 _17968__1483/HI net1483 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_95_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13344__A1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11254_ _06906_ _07081_ _07084_ _05263_ _06903_ vssd1 vssd1 vccd1 vccd1 _07594_ sky130_fd_sc_hd__o221a_1
X_14042_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[3\] _04265_ _04267_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[27\]
+ _04330_ vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__a221o_1
XANTENNA__10158__A1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10704__B net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10205_ net1140 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[8\] net968 vssd1
+ vssd1 vccd1 vccd1 _06545_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_52_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11185_ _07375_ _07523_ _07524_ net338 vssd1 vssd1 vccd1 vccd1 _07525_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17801_ clknet_leaf_121_wb_clk_i net2713 _01741_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[71\]
+ sky130_fd_sc_hd__dfrtp_1
X_10136_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[11\] net819 net804 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06476_ sky130_fd_sc_hd__a22o_1
X_15993_ net1410 vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__inv_2
XANTENNA__13647__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17732_ clknet_leaf_125_wb_clk_i _03408_ _01672_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11658__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10067_ _06280_ _06283_ vssd1 vssd1 vccd1 vccd1 _06407_ sky130_fd_sc_hd__or2_1
X_14944_ net1235 vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__inv_2
XANTENNA__12411__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08828__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09720__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16942__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17663_ clknet_leaf_3_wb_clk_i _03348_ _01604_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14875_ net1254 vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__inv_2
XANTENNA_clkload1_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16614_ clknet_leaf_73_wb_clk_i _02301_ _00597_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13826_ net2132 net831 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[19\]
+ sky130_fd_sc_hd__and2_1
X_17594_ clknet_leaf_89_wb_clk_i _03281_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10881__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14072__A2 _04258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16545_ clknet_leaf_6_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[11\]
+ _00528_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13757_ _04141_ _04142_ _04145_ vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__and3_2
XANTENNA__13280__B1 _04621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13846__A_N net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10969_ _06255_ _06410_ _07291_ vssd1 vssd1 vccd1 vccd1 _07309_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10094__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12708_ net2522 net227 net383 vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__mux2_1
X_16476_ clknet_leaf_151_wb_clk_i _02230_ _00459_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13688_ team_01_WB.instance_to_wrap.cpu.c0.count\[15\] _04109_ vssd1 vssd1 vccd1
+ vccd1 _04111_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08563__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15427_ net1221 vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__inv_2
X_12639_ net2976 net259 net393 vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13583__A1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09956__A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15358_ net1345 vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__inv_2
XANTENNA__09251__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold205 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[21\] vssd1 vssd1 vccd1 vccd1
+ net1740 sky130_fd_sc_hd__dlygate4sd3_1
X_14309_ net1324 vssd1 vssd1 vccd1 vccd1 _00103_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold216 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1751 sky130_fd_sc_hd__dlygate4sd3_1
X_15289_ net1238 vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__inv_2
Xhold227 team_01_WB.instance_to_wrap.a1.ADR_I\[9\] vssd1 vssd1 vccd1 vccd1 net1762
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 team_01_WB.instance_to_wrap.a1.ADR_I\[12\] vssd1 vssd1 vccd1 vccd1 net1773
+ sky130_fd_sc_hd__dlygate4sd3_1
X_17028_ clknet_leaf_84_wb_clk_i _02715_ _01011_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_113_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold249 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1784 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout707 net708 vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__clkbuf_4
X_09850_ net376 net342 _05416_ net560 vssd1 vssd1 vccd1 vccd1 _06190_ sky130_fd_sc_hd__a31o_1
XANTENNA__11897__A1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout718 net719 vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__clkbuf_4
X_08801_ net1093 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[0\] net917 vssd1
+ vssd1 vccd1 vccd1 _05141_ sky130_fd_sc_hd__and3_1
XANTENNA__17681__Q team_01_WB.instance_to_wrap.cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09781_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[15\] net737 net731 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12321__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08732_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[5\] net663 _05048_ _05050_
+ _05055_ vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_0_Left_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10630__A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09711__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08663_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[10\] net656 _04982_
+ _04984_ _04992_ vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08738__C net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08594_ net1104 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[15\] net909
+ net692 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[15\] vssd1 vssd1 vccd1
+ vccd1 _04934_ sky130_fd_sc_hd__a32o_1
XFILLER_0_89_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14063__A2 _04254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08278__A0 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13271__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_138_Right_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout340_A _06495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1082_A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10085__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09569__C net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09490__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09215_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[17\] net684 _05534_
+ _05537_ _05550_ vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_146_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12991__S net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09146_ _05482_ _05483_ _05484_ _05485_ vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_20_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13388__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09077_ _05416_ vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1135_X net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_49_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08028_ team_01_WB.instance_to_wrap.cpu.K0.keyvalid _04523_ vssd1 vssd1 vccd1 vccd1
+ _04524_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_9_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold750 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2285 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout974_A _04640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold761 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2296 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold772 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[18\] vssd1 vssd1 vccd1 vccd1
+ net2307 sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2318 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1302_X net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold794 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2329 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13835__B net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09979_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[2\] net787 net780 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06319_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout762_X net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13629__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12231__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12990_ net2609 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[104\] net852 vssd1 vssd1
+ vccd1 vccd1 _02135_ sky130_fd_sc_hd__mux2_1
Xhold1450 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2985 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08648__C net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1461 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 net2996
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1472 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net3007 sky130_fd_sc_hd__dlygate4sd3_1
X_11941_ net1943 net263 net476 vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__mux2_1
XANTENNA__14039__C1 net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13869__A_N net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1483 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net3018 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1494 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net3029 sky130_fd_sc_hd__dlygate4sd3_1
X_14660_ net1307 vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__inv_2
X_11872_ net2365 net238 net483 vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13611_ _03897_ _04051_ _03891_ vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__a21oi_1
X_10823_ _07055_ _07161_ vssd1 vssd1 vccd1 vccd1 _07163_ sky130_fd_sc_hd__nor2_1
XANTENNA__08808__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14591_ net1402 vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16330_ clknet_leaf_101_wb_clk_i _02084_ _00313_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[53\]
+ sky130_fd_sc_hd__dfstp_1
X_13542_ net185 _03993_ _03994_ net723 vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__a211o_1
XFILLER_0_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10754_ _04844_ net510 vssd1 vssd1 vccd1 vccd1 _07094_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_45_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09481__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16261_ clknet_leaf_151_wb_clk_i net1676 _00249_ vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13473_ _03855_ _03921_ _03933_ _03853_ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__o211a_1
X_10685_ net514 _07023_ _07024_ vssd1 vssd1 vccd1 vccd1 _07025_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_97_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18000_ net635 vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__clkbuf_1
X_15212_ net1259 vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13565__A1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10418__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09769__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12424_ net2914 net188 net415 vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16192_ clknet_leaf_1_wb_clk_i _01952_ _00180_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09233__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15143_ net1390 vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12406__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12355_ net2696 net315 net429 vssd1 vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13317__A1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11306_ _07645_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] _07638_ vssd1
+ vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__mux2_1
X_12286_ net2377 net309 net436 vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15074_ net1351 vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14025_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[10\] _04226_ _04251_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[82\]
+ _04314_ vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__a221o_1
X_11237_ net523 _07219_ _07576_ vssd1 vssd1 vccd1 vccd1 _07577_ sky130_fd_sc_hd__o21a_1
X_11168_ _07323_ _07438_ _07491_ _07507_ vssd1 vssd1 vccd1 vccd1 _07508_ sky130_fd_sc_hd__and4bb_1
XANTENNA__10551__A1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08398__Y _04738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10119_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[6\] net805 net758 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06459_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12141__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11099_ _06406_ _06408_ vssd1 vssd1 vccd1 vccd1 _07439_ sky130_fd_sc_hd__and2_1
X_15976_ net1354 vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17715_ clknet_leaf_115_wb_clk_i _03399_ _01656_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08558__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14927_ net1385 vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11980__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17646_ clknet_leaf_150_wb_clk_i _03331_ _01587_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14858_ net1374 vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__inv_2
XANTENNA__08855__A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14045__A2 _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13809_ net2996 net832 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[2\]
+ sky130_fd_sc_hd__and2_1
X_17577_ clknet_leaf_94_wb_clk_i _03264_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14789_ net1262 vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16528_ clknet_leaf_159_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[26\]
+ _00511_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16459_ clknet_leaf_28_wb_clk_i _02213_ _00442_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09000_ net1100 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[9\] net936 vssd1
+ vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__and3_1
XFILLER_0_73_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09224__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17676__Q team_01_WB.instance_to_wrap.cpu.DM0.readdata\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12316__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10790__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09902_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[5\] _04654_ net775 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06242_ sky130_fd_sc_hd__a22o_1
Xfanout504 _06779_ vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__buf_2
Xfanout515 net516 vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__clkbuf_4
Xfanout526 net527 vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__dlymetal6s2s_1
X_09833_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[13\] net821 net797 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06173_ sky130_fd_sc_hd__a22o_1
Xfanout537 net538 vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__clkbuf_2
Xfanout548 net549 vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10542__A1 _06881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout559 net560 vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout388_A _03569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10998__C _06902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12051__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09764_ _06068_ _06069_ vssd1 vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__or2_1
X_08715_ net1018 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[5\] net936 vssd1
+ vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__and3_1
X_09695_ net509 _06033_ vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__nor2_1
XANTENNA__13492__B1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11890__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout555_A net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_99_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08646_ net1020 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[10\] net916
+ vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17967__1482 vssd1 vssd1 vccd1 vccd1 _17967__1482/HI net1482 sky130_fd_sc_hd__conb_1
XANTENNA__14036__A2 _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13390__B _05705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout343_X net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08577_ _04904_ _04908_ _04912_ _04916_ vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_25_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10058__B1 _06396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09999__B1 _06337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09299__C net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout510_X net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout608_X net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13547__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09596__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10470_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[26\] net766 net624 vssd1
+ vssd1 vccd1 vccd1 _06810_ sky130_fd_sc_hd__o21a_1
XANTENNA__09215__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08931__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09129_ net1104 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[14\] net880
+ vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__and3_1
XFILLER_0_150_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12226__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12140_ net2105 net262 net452 vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__mux2_1
XANTENNA__10781__A1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout977_X net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12071_ net1739 net237 net459 vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__mux2_1
Xhold580 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 net2115
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12750__A net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold591 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2126 sky130_fd_sc_hd__dlygate4sd3_1
X_11022_ _05529_ net371 vssd1 vssd1 vccd1 vccd1 _07362_ sky130_fd_sc_hd__nand2_1
X_15830_ net1339 vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15761_ net1198 vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12973_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[113\] net1800 net866 vssd1 vssd1
+ vccd1 vccd1 _02152_ sky130_fd_sc_hd__mux2_1
X_17500_ clknet_leaf_58_wb_clk_i _03187_ _01483_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1280 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[89\] vssd1 vssd1 vccd1 vccd1
+ net2815 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09151__A1 _05490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1291 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2826 sky130_fd_sc_hd__dlygate4sd3_1
X_14712_ net1191 vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__inv_2
X_11924_ net2173 net290 net480 vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15692_ net1260 vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14027__A2 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17431_ clknet_leaf_13_wb_clk_i _03118_ _01414_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_14643_ net1256 vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__inv_2
X_11855_ net2734 net305 net490 vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_72_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10049__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10806_ _07144_ _07145_ _07142_ vssd1 vssd1 vccd1 vccd1 _07146_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17362_ clknet_leaf_144_wb_clk_i _03049_ _01345_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14574_ net1401 vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__inv_2
X_11786_ net2059 net311 net497 vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09454__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_25 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16313_ clknet_leaf_118_wb_clk_i _02067_ _00296_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[36\]
+ sky130_fd_sc_hd__dfstp_1
X_13525_ net988 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] _03979_ _03980_
+ vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09002__C net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10737_ _06966_ _06967_ _06964_ vssd1 vssd1 vccd1 vccd1 _07077_ sky130_fd_sc_hd__a21oi_1
X_17293_ clknet_leaf_68_wb_clk_i _02980_ _01276_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16244_ clknet_leaf_140_wb_clk_i net1654 _00232_ vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__dfrtp_1
X_13456_ _03914_ _03916_ vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__and2_1
XFILLER_0_153_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_153_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10668_ net547 net372 _07007_ vssd1 vssd1 vccd1 vccd1 _07008_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_152_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10716__Y _07056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12407_ net3168 net231 net421 vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16175_ clknet_leaf_6_wb_clk_i _01935_ _00163_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12136__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13387_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] _05727_ vssd1 vssd1
+ vccd1 vccd1 _03848_ sky130_fd_sc_hd__and2_1
X_10599_ net550 _06562_ vssd1 vssd1 vccd1 vccd1 _06939_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__buf_2
X_15126_ net1246 vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__inv_2
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__buf_2
Xoutput129 net129 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__buf_2
X_12338_ net2050 net234 net427 vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_110_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_81_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11975__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15057_ net1393 vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__inv_2
X_12269_ net2614 net244 net437 vssd1 vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__mux2_1
X_14008_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[57\] _04258_ _04264_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[105\]
+ _04298_ vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__a221o_1
XANTENNA__09672__C net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_133_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11721__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11276__A _06919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09390__A1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17636__CLK clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15959_ net1412 vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_108_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12816__A3 _03639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08500_ _04717_ _04752_ _04838_ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__or3_1
XANTENNA__10288__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09480_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[30\] net693 net662 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_90_Left_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08585__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08431_ net1025 net924 vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__and2_2
XANTENNA__16575__Q team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17629_ clknet_leaf_3_wb_clk_i _03314_ _01570_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08362_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[30\] net742 _04681_
+ _04677_ _04670_ vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_18_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08293_ net1161 net1164 net1166 net1158 vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_15_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13529__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10460__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08751__C net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1030 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12046__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout303_A _07912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1045_A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10212__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10763__A1 _06958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11885__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1212_A net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout301 net303 vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__buf_2
Xfanout312 _07931_ vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__buf_1
XANTENNA__09905__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout323 net326 vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__buf_2
Xfanout334 _06918_ vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout672_A _04794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout345 net347 vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__buf_2
XANTENNA__10802__B net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08479__B net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13953__X _04245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout356 _03655_ vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09381__A1 net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09816_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[14\] net766 vssd1 vssd1
+ vccd1 vccd1 _06156_ sky130_fd_sc_hd__or2_1
Xfanout367 _07759_ vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout389 _03569_ vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__buf_6
XANTENNA__10521__C net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_129_Left_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12268__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09747_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[20\] net742 _06072_
+ _06075_ _06076_ vssd1 vssd1 vccd1 vccd1 _06087_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout460_X net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout937_A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout558_X net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09678_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[22\] net815 net777 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__a22o_1
XANTENNA__14009__A2 _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08926__C net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08629_ net601 _04968_ _04949_ vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_139_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout725_X net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11640_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] _07817_ vssd1 vssd1
+ vccd1 vccd1 _07850_ sky130_fd_sc_hd__xor2_1
XFILLER_0_65_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09436__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11243__A2 _07527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11571_ net3085 net152 team_01_WB.instance_to_wrap.cpu.K0.next_state vssd1 vssd1
+ vccd1 vccd1 _03271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_64_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13310_ team_01_WB.instance_to_wrap.cpu.f0.i\[20\] _07707_ vssd1 vssd1 vccd1 vccd1
+ _03792_ sky130_fd_sc_hd__or2_1
X_10522_ net1080 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[31\] net891
+ vssd1 vssd1 vccd1 vccd1 _06862_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_138_Left_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14290_ net1346 vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13241_ net2907 net354 net350 team_01_WB.instance_to_wrap.cpu.f0.i\[9\] vssd1 vssd1
+ vccd1 vccd1 _01909_ sky130_fd_sc_hd__a22o_1
X_10453_ net1147 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[26\] net957
+ vssd1 vssd1 vccd1 vccd1 _06793_ sky130_fd_sc_hd__and3_1
XFILLER_0_150_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12743__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10384_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[16\] net818 net781 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06724_ sky130_fd_sc_hd__a22o_1
XANTENNA_input66_A wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13172_ net134 net848 net840 net1656 vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__a22o_1
XANTENNA__11795__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12123_ net2117 net290 net456 vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__mux2_1
X_17980_ net1495 vssd1 vssd1 vccd1 vccd1 la_data_out[22] sky130_fd_sc_hd__buf_2
X_12054_ net2018 net307 net466 vssd1 vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__mux2_1
XANTENNA__16533__CLK clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16931_ clknet_leaf_25_wb_clk_i _02618_ _00914_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11005_ _05729_ _06812_ vssd1 vssd1 vccd1 vccd1 _07345_ sky130_fd_sc_hd__and2_1
X_16862_ clknet_leaf_80_wb_clk_i _02549_ _00845_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout890 _04799_ vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__buf_4
X_15813_ net1200 vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__inv_2
X_16793_ clknet_leaf_103_wb_clk_i _02480_ _00776_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15744_ net1232 vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12956_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[4\] _05110_ net1038 vssd1
+ vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11907_ net2590 net267 net480 vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__mux2_1
X_15675_ net1255 vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[26\] _03665_ net1037 vssd1
+ vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17414_ clknet_leaf_103_wb_clk_i _03101_ _01397_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14626_ net1262 vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09788__X _06128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11838_ net1944 net271 net489 vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_155_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09427__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17345_ clknet_leaf_50_wb_clk_i _03032_ _01328_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14557_ net1410 vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__inv_2
X_11769_ net1912 net243 net496 vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13508_ net724 _07056_ net987 vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__a21oi_1
X_17276_ clknet_leaf_59_wb_clk_i _02963_ _01259_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14488_ net1347 vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__inv_2
XANTENNA__09667__C net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_0__f_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_0__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__08571__C net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16227_ clknet_leaf_133_wb_clk_i net1707 _00215_ vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__dfrtp_1
X_13439_ _03883_ _03896_ _03899_ vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__o21a_1
XFILLER_0_140_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16158_ clknet_leaf_134_wb_clk_i _01921_ _00146_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10745__A1 _06906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17966__1481 vssd1 vssd1 vccd1 vccd1 _17966__1481/HI net1481 sky130_fd_sc_hd__conb_1
XFILLER_0_122_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15109_ net1262 vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__inv_2
X_08980_ _05307_ _05311_ net619 _05319_ vssd1 vssd1 vccd1 vccd1 _05320_ sky130_fd_sc_hd__and4bb_1
X_16089_ clknet_leaf_132_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[11\]
+ _00077_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08299__B net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10341__C net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09601_ net1146 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[24\] net957
+ vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_127_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09532_ net1152 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[28\] net979
+ vssd1 vssd1 vccd1 vccd1 _05872_ sky130_fd_sc_hd__and3_1
XANTENNA__08746__C net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09463_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] net710 net594 vssd1 vssd1
+ vccd1 vccd1 _05803_ sky130_fd_sc_hd__a21o_2
XANTENNA__08874__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout253_A net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10681__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08414_ net711 _04751_ _04752_ vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__nor3_2
XFILLER_0_59_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09394_ net559 _05659_ vssd1 vssd1 vccd1 vccd1 _05734_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08345_ net991 net958 vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08626__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout420_A net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1162_A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout518_A _05260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08276_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[5\] net2036 net1042 vssd1 vssd1
+ vccd1 vccd1 _03411_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13948__X _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1427_A net1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout887_A _04799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12504__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1107 net1114 vssd1 vssd1 vccd1 vccd1 net1107 sky130_fd_sc_hd__clkbuf_2
Xfanout1118 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[23\] vssd1 vssd1 vccd1 vccd1
+ net1118 sky130_fd_sc_hd__buf_2
XFILLER_0_100_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout675_X net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1129 net1130 vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13150__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_111_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_111_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_156_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout186 _07639_ vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__clkbuf_4
Xfanout197 _07633_ vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__buf_2
XANTENNA__13843__B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout842_X net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12810_ net1714 net640 net608 _03635_ vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__a22o_1
X_13790_ net1184 _04160_ vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_83_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[28\] _07088_ net1034 vssd1 vssd1
+ vccd1 vccd1 _03588_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15460_ net1219 vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__inv_2
X_12672_ net3065 net259 net389 vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ net1359 vssd1 vssd1 vccd1 vccd1 _00205_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_146_Left_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11623_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[27\] _07566_ net715 vssd1 vssd1
+ vccd1 vccd1 _07836_ sky130_fd_sc_hd__mux2_1
X_15391_ net1318 vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__inv_2
XANTENNA__08617__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17130_ clknet_leaf_10_wb_clk_i _02817_ _01113_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_14342_ net1338 vssd1 vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__inv_2
X_11554_ net37 net36 net35 net34 vssd1 vssd1 vccd1 vccd1 _07786_ sky130_fd_sc_hd__nor4_1
X_17061_ clknet_leaf_52_wb_clk_i _02748_ _01044_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10505_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[31\] net759 net754 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06845_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14273_ net1340 vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11485_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[20\] net580 vssd1 vssd1 vccd1
+ vccd1 _07770_ sky130_fd_sc_hd__nand2_1
X_16012_ net1348 vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13224_ net3040 net353 net349 team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1
+ vccd1 vccd1 _01926_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10436_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[27\] net739 _06774_ _06775_
+ net768 vssd1 vssd1 vccd1 vccd1 _06776_ sky130_fd_sc_hd__a2111o_1
XANTENNA_input69_X net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13155_ net1706 net850 net842 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[21\] vssd1
+ vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__a22o_1
XANTENNA__12414__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10367_ net581 _06706_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] net625
+ vssd1 vssd1 vccd1 vccd1 _06707_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_27_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12106_ net1752 net267 net456 vssd1 vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_155_Left_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10298_ net559 _04919_ _05731_ _06637_ vssd1 vssd1 vccd1 vccd1 _06638_ sky130_fd_sc_hd__a22oi_2
X_13086_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[0\] net3069 net852 vssd1 vssd1
+ vccd1 vccd1 _02039_ sky130_fd_sc_hd__mux2_1
X_17963_ net1478 vssd1 vssd1 vccd1 vccd1 la_data_out[5] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_148_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12037_ net2494 net270 net463 vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__mux2_1
X_16914_ clknet_leaf_143_wb_clk_i _02601_ _00897_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17894_ net1516 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
XANTENNA__09896__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09950__C _04660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16845_ clknet_leaf_68_wb_clk_i _02532_ _00828_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_144_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16776_ clknet_leaf_63_wb_clk_i _02463_ _00759_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13988_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[88\] _04241_ _04250_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[120\]
+ _04270_ vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__a221o_1
XANTENNA__09648__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08566__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15727_ net1300 vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_122_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08856__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12939_ net1798 net870 net357 _03702_ vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15658_ net1377 vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__inv_2
XANTENNA__08863__A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14609_ net1340 vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15589_ net1263 vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08130_ team_01_WB.instance_to_wrap.cpu.f0.i\[30\] _04493_ team_01_WB.instance_to_wrap.cpu.f0.num\[7\]
+ _04486_ _04582_ vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__a221o_1
XFILLER_0_56_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17328_ clknet_leaf_146_wb_clk_i _03015_ _01311_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08061_ _04522_ _04528_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17259_ clknet_leaf_8_wb_clk_i _02946_ _01242_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09694__A net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17684__Q team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_113_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08387__A2 _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10194__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08963_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\] net596 vssd1 vssd1 vccd1
+ vccd1 _05303_ sky130_fd_sc_hd__nand2_1
XANTENNA__13132__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08894_ net1025 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[2\] net931 vssd1
+ vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__and3_1
XANTENNA__10071__C net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1008_A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout468_A net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14093__B1 _04265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09515_ _05851_ _05852_ _05853_ _05854_ vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__or4_1
XANTENNA__08476__C net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout256_X net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1377_A net1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10654__A0 _05898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09446_ net1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[29\] net920 vssd1
+ vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08773__A net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17859__Q team_01_WB.instance_to_wrap.cpu.f0.read_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_47_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout802_A _04643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10367__X _06707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout423_X net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09377_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[26\] _04808_ net649
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[26\] _05714_ vssd1 vssd1 vccd1
+ vccd1 _05717_ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12946__A2 _07757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08328_ net1130 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[30\] net975
+ vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__and3_1
XFILLER_0_145_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10957__A1 _06919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09811__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09100__C net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08259_ net3033 net3186 net1042 vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1332_X net1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13838__B net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11270_ _07605_ _07608_ _07609_ vssd1 vssd1 vccd1 vccd1 _07610_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout792_X net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10814__Y _07154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10221_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[8\] net763 net622 vssd1
+ vssd1 vccd1 vccd1 _06561_ sky130_fd_sc_hd__o21a_1
XANTENNA__12234__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10543__A net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10152_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[11\] net742 net734 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[11\]
+ _06491_ vssd1 vssd1 vccd1 vccd1 _06492_ sky130_fd_sc_hd__a221o_1
XANTENNA__08013__A net1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13659__B1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13123__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10083_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[7\] net772 net744 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[7\]
+ _06416_ vssd1 vssd1 vccd1 vccd1 _06423_ sky130_fd_sc_hd__a221o_1
XANTENNA__10830__X _07170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14960_ net1272 vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_7_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold9 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[1\] vssd1 vssd1 vccd1 vccd1
+ net1544 sky130_fd_sc_hd__dlygate4sd3_1
X_13911_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[9\] _04207_ vssd1 vssd1 vccd1
+ vccd1 _04209_ sky130_fd_sc_hd__and2_1
X_14891_ net1397 vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__inv_2
XANTENNA_input29_A DAT_I[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08300__X _04640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16630_ clknet_leaf_30_wb_clk_i _02317_ _00613_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10893__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13842_ net1179 net1066 net3172 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[3\]
+ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_18_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14084__B1 _04259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16561_ clknet_leaf_159_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[27\]
+ _00544_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13773_ _04154_ _04158_ vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__nor2_1
XANTENNA__12634__A1 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10985_ net547 _06398_ vssd1 vssd1 vccd1 vccd1 _07325_ sky130_fd_sc_hd__nor2_1
XANTENNA__10645__A0 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15512_ net1214 vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12724_ net1032 _03573_ _03574_ net1175 vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__a211o_1
XFILLER_0_29_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17965__1480 vssd1 vssd1 vccd1 vccd1 _17965__1480/HI net1480 sky130_fd_sc_hd__conb_1
X_16492_ clknet_leaf_151_wb_clk_i _02246_ _00475_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12917__B net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15443_ net1419 vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__inv_2
X_12655_ net2855 net188 net387 vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__mux2_1
XANTENNA__12409__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11606_ _07796_ _07822_ net611 vssd1 vssd1 vccd1 vccd1 _07823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15374_ net1292 vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12586_ net2787 net314 net402 vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__mux2_1
XANTENNA__09263__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09802__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17113_ clknet_leaf_104_wb_clk_i _02800_ _01096_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11070__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14325_ net1331 vssd1 vssd1 vccd1 vccd1 _00119_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11537_ net2556 net1174 net589 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[16\] vssd1
+ vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__a22o_1
XANTENNA__09010__C net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold409 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1944 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_78_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17044_ clknet_leaf_22_wb_clk_i _02731_ _01027_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_14256_ net1226 vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__inv_2
X_11468_ net366 _07761_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[29\] net874
+ vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_123_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13207_ net32 net838 _03738_ net3157 vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__a22o_1
X_10419_ net1133 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[27\] net957
+ vssd1 vssd1 vccd1 vccd1 _06759_ sky130_fd_sc_hd__and3b_1
X_14187_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[13\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[12\]
+ _04453_ vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__and3_1
XANTENNA__12144__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10176__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11399_ team_01_WB.instance_to_wrap.cpu.f0.i\[25\] _07695_ vssd1 vssd1 vccd1 vccd1
+ _07723_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_74_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ net1651 net846 net634 team_01_WB.instance_to_wrap.a1.ADR_I\[5\] vssd1 vssd1
+ vccd1 vccd1 _02003_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_146_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11983__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13114__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17946_ net1461 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
X_13069_ net2238 net2205 net865 vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__mux2_1
Xhold1109 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2644 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09869__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08858__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17877_ clknet_leaf_139_wb_clk_i _03552_ _01817_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11284__A _07135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16828_ clknet_leaf_57_wb_clk_i _02515_ _00811_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14075__B1 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16759_ clknet_leaf_15_wb_clk_i _02446_ _00742_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_09300_ net1084 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[22\] net879
+ vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__and3_1
XANTENNA__10636__A0 _06912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17679__Q team_01_WB.instance_to_wrap.cpu.f0.i\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_152_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09231_ net1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[21\] net890 vssd1
+ vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__and3_1
XANTENNA__12319__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12928__A2 _07757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09162_ net1091 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[16\] net930
+ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__and3_1
XANTENNA__08057__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09254__B1 _05593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08880__X _05220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08113_ team_01_WB.instance_to_wrap.cpu.f0.i\[29\] team_01_WB.instance_to_wrap.cpu.f0.num\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__xor2_1
XFILLER_0_146_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13939__A team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09093_ net1013 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[13\] net922 vssd1
+ vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout216_A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08044_ net1591 net570 net346 team_01_WB.instance_to_wrap.cpu.f0.i\[11\] vssd1 vssd1
+ vccd1 vccd1 _03547_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold910 _02088_ vssd1 vssd1 vccd1 vccd1 net2445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2456 sky130_fd_sc_hd__dlygate4sd3_1
Xhold932 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[14\] vssd1 vssd1 vccd1 vccd1 net2467
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_80 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold943 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2478 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12054__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold954 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2489 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10167__A2 _04667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold965 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2500 sky130_fd_sc_hd__dlygate4sd3_1
Xhold976 team_01_WB.instance_to_wrap.cpu.f0.num\[0\] vssd1 vssd1 vccd1 vccd1 net2511
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2522 sky130_fd_sc_hd__dlygate4sd3_1
X_17989__1504 vssd1 vssd1 vccd1 vccd1 _17989__1504/HI net1504 sky130_fd_sc_hd__conb_1
Xhold998 _02146_ vssd1 vssd1 vccd1 vccd1 net2533 sky130_fd_sc_hd__dlygate4sd3_1
X_09995_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[2\] net775 net737 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06335_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13096__D net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11893__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11746__X _07935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08780__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08946_ net1028 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[6\] net894 vssd1
+ vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_32_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1610 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net3145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1621 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net3156 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1632 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net3167 sky130_fd_sc_hd__dlygate4sd3_1
X_08877_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[3\] net675 net660 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[3\]
+ net706 vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout752_A _04678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1643 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 net3178
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10810__B net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout373_X net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13961__X _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08532__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10088__D1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09599__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10770_ _07103_ _07109_ vssd1 vssd1 vccd1 vccd1 _07110_ sky130_fd_sc_hd__or2_1
XANTENNA__08934__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09429_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[28\] net667 net665 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[28\]
+ _05768_ vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__a221o_1
XANTENNA__12229__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout805_X net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12440_ net2371 net229 net417 vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08599__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13592__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12371_ net1808 net236 net423 vssd1 vssd1 vccd1 vccd1 _02625_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14110_ _04217_ _04231_ _04239_ vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__and3_1
X_11322_ _07657_ net2109 _07655_ vssd1 vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__mux2_1
X_15090_ net1266 vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_95_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14041_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[75\] _04268_ _04289_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__a22o_1
X_11253_ _07055_ _07278_ vssd1 vssd1 vccd1 vccd1 _07593_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10204_ net1139 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[8\] net945 vssd1
+ vssd1 vccd1 vccd1 _06544_ sky130_fd_sc_hd__and3_1
X_11184_ _07014_ _07149_ _07242_ net522 vssd1 vssd1 vccd1 vccd1 _07524_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17800_ clknet_leaf_117_wb_clk_i net2724 _01740_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[70\]
+ sky130_fd_sc_hd__dfrtp_1
X_10135_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[11\] net791 net752 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[11\]
+ _06473_ vssd1 vssd1 vccd1 vccd1 _06475_ sky130_fd_sc_hd__a221o_1
X_15992_ net1364 vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__inv_2
XANTENNA__13501__C1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10066_ _06404_ _06405_ _06316_ vssd1 vssd1 vccd1 vccd1 _06406_ sky130_fd_sc_hd__a21oi_2
X_14943_ net1317 vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__inv_2
X_17731_ clknet_leaf_125_wb_clk_i _03407_ _01671_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11658__A2 _07171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17662_ clknet_leaf_0_wb_clk_i _03347_ _01603_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_14874_ net1371 vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__inv_2
X_16613_ clknet_leaf_51_wb_clk_i _02300_ _00596_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13825_ net2055 net830 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[18\]
+ sky130_fd_sc_hd__and2_1
X_17593_ clknet_leaf_89_wb_clk_i _03280_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09005__C net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16544_ clknet_leaf_6_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[10\]
+ _00527_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13756_ _04143_ _04144_ vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__nor2_1
X_10968_ _07276_ _07306_ _07307_ _07299_ vssd1 vssd1 vccd1 vccd1 _07308_ sky130_fd_sc_hd__o211a_2
XFILLER_0_156_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12707_ net2835 net284 net386 vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__mux2_1
XANTENNA__09302__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11291__B1 _06960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16475_ clknet_leaf_140_wb_clk_i _02229_ _00458_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12139__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13687_ team_01_WB.instance_to_wrap.cpu.c0.count\[15\] _04109_ vssd1 vssd1 vccd1
+ vccd1 _04110_ sky130_fd_sc_hd__or2_1
X_10899_ net557 _07238_ _06963_ vssd1 vssd1 vccd1 vccd1 _07239_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_139_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15426_ net1319 vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__inv_2
XANTENNA__08039__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12638_ net2777 net229 net392 vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11978__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13583__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15357_ net1315 vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12569_ net2037 net234 net399 vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_117_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10397__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14308_ net1324 vssd1 vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__inv_2
XANTENNA__12791__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15288_ net1215 vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__inv_2
Xhold206 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1741 sky130_fd_sc_hd__dlygate4sd3_1
Xhold217 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1752 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09675__C net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold228 team_01_WB.instance_to_wrap.cpu.f0.write_data\[6\] vssd1 vssd1 vccd1 vccd1
+ net1763 sky130_fd_sc_hd__dlygate4sd3_1
X_17027_ clknet_leaf_23_wb_clk_i _02714_ _01010_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_113_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold239 net99 vssd1 vssd1 vccd1 vccd1 net1774 sky130_fd_sc_hd__dlygate4sd3_1
X_14239_ net1206 vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__inv_2
XANTENNA__16617__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10149__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout708 _04757_ vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__buf_4
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout719 _04722_ vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__buf_2
X_08800_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[0\] net662 _05138_ _05139_
+ net705 vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08762__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09780_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[15\] net757 net735 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__a22o_1
XANTENNA__12602__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08731_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[5\] net688 _05057_ _05058_
+ _05063_ vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__a2111o_1
X_17929_ net1446 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
XANTENNA__12846__A1 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10630__B net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1290 net1292 vssd1 vssd1 vccd1 vccd1 net1290 sky130_fd_sc_hd__buf_4
XANTENNA__10857__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_89_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08662_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[10\] net694 _04973_
+ _04976_ net706 vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__a2111o_1
XANTENNA__14048__B1 _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08593_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[15\] net652 _04921_
+ _04924_ _04927_ vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_152_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10609__A0 _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08754__C net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09212__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12049__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout333_A net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1075_A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09214_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[17\] net687 _05541_ _05546_
+ _05551_ vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13559__C1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11888__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09145_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[14\] net673 _05470_ _05474_
+ _05478_ vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_101_Left_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout500_A net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1242_A net1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10388__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09242__A3 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12782__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09076_ _05380_ _05415_ net603 vssd1 vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__mux2_2
XFILLER_0_32_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08027_ _04512_ _04522_ vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_9_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold740 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2275 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1030_X net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold751 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2286 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11337__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold762 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold773 _02057_ vssd1 vssd1 vccd1 vccd1 net2308 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09882__A net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold784 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2319 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout490_X net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold795 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2330 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11168__B_N _07438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_89_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_90_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12512__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09978_ net998 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[2\] net960 vssd1
+ vssd1 vccd1 vccd1 _06318_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_18_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08929_ net1111 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[6\] net890 vssd1
+ vssd1 vccd1 vccd1 _05269_ sky130_fd_sc_hd__and3_1
XANTENNA__08929__C net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_110_Left_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout755_X net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1440 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2975 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1451 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2986 sky130_fd_sc_hd__dlygate4sd3_1
X_11940_ net2317 net268 net475 vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__mux2_1
XANTENNA__10848__B1 _07187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1462 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2997 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10312__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1473 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net3008 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1484 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[73\] vssd1 vssd1 vccd1 vccd1
+ net3019 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1495 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net3030 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13851__B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11871_ net2690 net270 net485 vssd1 vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout922_X net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13610_ _03883_ _03895_ vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__or2_1
X_10822_ net553 _07160_ _07161_ _06964_ vssd1 vssd1 vccd1 vccd1 _07162_ sky130_fd_sc_hd__a31o_1
XANTENNA__08269__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14590_ net1401 vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09122__A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13541_ net196 net192 _07854_ net642 vssd1 vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__o211a_1
XANTENNA__11371__B team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_95_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10753_ _06034_ _07091_ _06001_ vssd1 vssd1 vccd1 vccd1 _07093_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16260_ clknet_leaf_156_wb_clk_i net1692 _00248_ vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08383__D _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13472_ _03924_ _03929_ _03932_ vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__and3_1
XFILLER_0_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10684_ net537 _07022_ _06970_ vssd1 vssd1 vccd1 vccd1 _07024_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_97_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15211_ net1425 vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__inv_2
XANTENNA__11798__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12423_ _07942_ _07946_ net573 vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__and3_4
XFILLER_0_118_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13565__A2 _07135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16191_ clknet_leaf_1_wb_clk_i _01951_ _00179_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10379__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12773__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15142_ net1404 vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__inv_2
X_12354_ net2266 net318 net430 vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10715__B _06928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11305_ net727 _07476_ net187 _07644_ vssd1 vssd1 vccd1 vccd1 _07645_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15073_ net1280 vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12285_ net1854 net294 net438 vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14024_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[74\] _04235_ _04267_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__a22o_1
XANTENNA__09792__A net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11236_ _06906_ _07027_ _07033_ _05263_ net338 vssd1 vssd1 vccd1 vccd1 _07576_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_71_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_123_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_120_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12422__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11167_ _07502_ _07506_ _07494_ vssd1 vssd1 vccd1 vccd1 _07507_ sky130_fd_sc_hd__and3b_2
XFILLER_0_101_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10118_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[6\] net813 net786 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[6\]
+ _06444_ vssd1 vssd1 vccd1 vccd1 _06458_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12828__B2 _03648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11098_ _07431_ _07437_ _07339_ vssd1 vssd1 vccd1 vccd1 _07438_ sky130_fd_sc_hd__o21ai_4
X_15975_ net1413 vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__inv_2
X_17714_ clknet_leaf_125_wb_clk_i _03398_ _01655_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14926_ net1297 vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__inv_2
X_10049_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[0\] net776 net745 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06389_ sky130_fd_sc_hd__a22o_1
XANTENNA__10303__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17645_ clknet_leaf_157_wb_clk_i _03330_ _01586_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_69_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14857_ net1294 vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_86_831 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13808_ net2542 net833 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[1\]
+ sky130_fd_sc_hd__and2_1
X_17576_ clknet_leaf_94_wb_clk_i _03263_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__dfxtp_1
X_14788_ net1230 vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__inv_2
XANTENNA__09457__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08574__C net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16527_ clknet_leaf_159_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[25\]
+ _00510_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13739_ net1700 _04524_ team_01_WB.instance_to_wrap.cpu.f0.next_lcd_en vssd1 vssd1
+ vccd1 vccd1 _00024_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17988__1503 vssd1 vssd1 vccd1 vccd1 _17988__1503/HI net1503 sky130_fd_sc_hd__conb_1
XFILLER_0_129_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16458_ clknet_leaf_109_wb_clk_i _02212_ _00441_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15409_ net1393 vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16389_ clknet_leaf_122_wb_clk_i net2711 _00372_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[112\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12764__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10625__B net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10344__C net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09901_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[5\] net780 net740 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06241_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout505 _06636_ vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__clkbuf_4
Xfanout516 _05261_ vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__buf_4
X_09832_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[13\] net807 net742 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[13\]
+ _06171_ vssd1 vssd1 vccd1 vccd1 _06172_ sky130_fd_sc_hd__a221o_1
Xfanout527 _05223_ vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__clkbuf_2
X_17944__1459 vssd1 vssd1 vccd1 vccd1 _17944__1459/HI net1459 sky130_fd_sc_hd__conb_1
Xfanout538 net542 vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12332__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout549 _05151_ vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08749__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09763_ _06000_ _06034_ vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__nand2_1
XANTENNA__08111__A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout283_A _07908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08714_ net1097 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[5\] net884 vssd1
+ vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__and3_1
XANTENNA__16101__Q team_01_WB.instance_to_wrap.cpu.f0.data_adr\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09694_ net509 _06033_ vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08645_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[10\] net916
+ vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout450_A _07958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1192_A net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08576_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[19\] net698 _04913_
+ _04914_ _04915_ vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09448__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13244__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_49_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08484__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09999__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_136_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_136_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout336_X net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout715_A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08781__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13399__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12507__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout503_X net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1245_X net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09128_ net1110 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[14\] net893
+ vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09620__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09059_ net1029 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[12\] net880
+ vssd1 vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__and3_1
XFILLER_0_130_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12070_ net2348 net271 net461 vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold570 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2105 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout872_X net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold581 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2116 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12750__B _07579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold592 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2127 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08726__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11021_ _07360_ vssd1 vssd1 vccd1 vccd1 _07361_ sky130_fd_sc_hd__inv_2
XANTENNA__12242__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10533__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11366__B team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_99_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15760_ net1342 vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__inv_2
X_12972_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[114\] net1742 net863 vssd1 vssd1
+ vccd1 vccd1 _02153_ sky130_fd_sc_hd__mux2_1
XANTENNA__09687__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1270 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2805 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input11_A DAT_I[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11923_ net3169 net314 net481 vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__mux2_1
X_14711_ net1191 vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__inv_2
Xhold1281 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[24\] vssd1 vssd1 vccd1 vccd1
+ net2816 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15691_ net1423 vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__inv_2
XANTENNA__11494__B1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1292 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2827 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_47_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14642_ net1282 vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__inv_2
X_17430_ clknet_leaf_30_wb_clk_i _03117_ _01413_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11854_ net2471 net312 net490 vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1036 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10805_ _05657_ net331 _07143_ net336 net369 vssd1 vssd1 vccd1 vccd1 _07145_ sky130_fd_sc_hd__a221o_1
X_17361_ clknet_leaf_113_wb_clk_i _03048_ _01344_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14573_ net1410 vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11785_ net1727 net293 net496 vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_136_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13524_ net721 _07588_ net1074 vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__o21a_1
X_16312_ clknet_leaf_97_wb_clk_i _02066_ _00295_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10736_ _07074_ _07075_ _07072_ vssd1 vssd1 vccd1 vccd1 _07076_ sky130_fd_sc_hd__o21ba_1
X_17292_ clknet_leaf_147_wb_clk_i _02979_ _01275_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16243_ clknet_leaf_141_wb_clk_i net1652 _00231_ vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13455_ _03859_ _03915_ vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__and2b_1
XFILLER_0_82_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10667_ net551 _06250_ vssd1 vssd1 vccd1 vccd1 _07007_ sky130_fd_sc_hd__nor2_1
XANTENNA__12417__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12406_ net2798 net261 net420 vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16174_ clknet_leaf_7_wb_clk_i _01934_ _00162_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09072__D1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13386_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] _05757_ vssd1 vssd1
+ vccd1 vccd1 _03847_ sky130_fd_sc_hd__and2_1
XANTENNA__09611__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10598_ _06936_ _06937_ net538 vssd1 vssd1 vccd1 vccd1 _06938_ sky130_fd_sc_hd__mux2_1
X_15125_ net1276 vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__inv_2
XANTENNA__10221__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[8\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__buf_2
X_12337_ net1934 net239 net427 vssd1 vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__mux2_1
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10164__C net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15056_ net1274 vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__inv_2
X_12268_ net2234 net202 net435 vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__mux2_1
X_14007_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[33\] _04230_ _04240_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[89\]
+ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11219_ _05758_ _07558_ vssd1 vssd1 vccd1 vccd1 _07559_ sky130_fd_sc_hd__nand2_1
XANTENNA__12152__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12199_ net1964 net204 net444 vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__mux2_1
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__buf_2
XANTENNA__10524__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08569__C net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11991__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15958_ net1407 vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_108_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13474__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09678__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08866__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13474__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09142__A2 _04789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09314__X _05654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14909_ net1241 vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15889_ net1401 vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08350__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08430_ net1119 net1123 net1126 net1117 vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__and4bb_4
XANTENNA__09033__Y _05373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17628_ clknet_leaf_3_wb_clk_i _03313_ _01569_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_53_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08361_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[30\] net819 net807 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17559_ clknet_leaf_17_wb_clk_i _03246_ _01542_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10339__C net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09697__A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08292_ net1139 net981 vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__and2_2
XFILLER_0_85_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09850__B1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16591__Q team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[23\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12327__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12737__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13859__A_N net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12752__A3 _03595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10923__X _07263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10074__C net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1038_A net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout302 net303 vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13162__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12062__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout313 net316 vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__buf_2
Xfanout324 net326 vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1205_A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout335 _06912_ vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__clkbuf_4
Xfanout346 net347 vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__clkbuf_2
X_09815_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[14\] net818 net762 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[14\]
+ _06154_ vssd1 vssd1 vccd1 vccd1 _06155_ sky130_fd_sc_hd__a221o_1
Xfanout357 net358 vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input3_A DAT_I[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout368 _06915_ vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__clkbuf_4
Xfanout379 net382 vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout665_A _04804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09746_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[20\] net811 _06074_ _06079_
+ _06082_ vssd1 vssd1 vccd1 vccd1 _06086_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09224__X _05564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11476__B1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09677_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[22\] net755 _06005_ _06007_
+ _06015_ vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout832_A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout453_X net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08628_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[11\] net701 _04961_ _04967_
+ vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__o22a_2
XTAP_TAPCELL_ROW_85_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09728__A_N net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08559_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[19\] net684 _04896_
+ _04897_ _04898_ vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_65_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout718_X net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10436__D1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11570_ team_01_WB.instance_to_wrap.cpu.K0.count\[1\] team_01_WB.instance_to_wrap.cpu.K0.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__or2_1
XFILLER_0_147_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09841__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08942__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10521_ net1003 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[31\] net940 vssd1
+ vssd1 vccd1 vccd1 _06861_ sky130_fd_sc_hd__and3_1
XANTENNA__12237__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13240_ net3058 net354 net350 team_01_WB.instance_to_wrap.cpu.f0.i\[10\] vssd1 vssd1
+ vccd1 vccd1 _01910_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_131_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10452_ net1148 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[26\] net971
+ vssd1 vssd1 vccd1 vccd1 _06792_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_131_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13171_ net1952 net848 net840 net1949 vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__a22o_1
X_10383_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[16\] net799 net787 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[16\]
+ _06722_ vssd1 vssd1 vccd1 vccd1 _06723_ sky130_fd_sc_hd__a221o_1
X_12122_ net1878 net313 net457 vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_33_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08303__X _04643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input59_A wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11377__A team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13153__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16930_ clknet_leaf_77_wb_clk_i _02617_ _00913_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12053_ net1822 net312 net466 vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__mux2_1
XANTENNA__11703__A1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10506__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17987__1502 vssd1 vssd1 vccd1 vccd1 _17987__1502/HI net1502 sky130_fd_sc_hd__conb_1
X_11004_ _07342_ _07343_ vssd1 vssd1 vccd1 vccd1 _07344_ sky130_fd_sc_hd__or2_1
XANTENNA__09372__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16861_ clknet_leaf_58_wb_clk_i _02548_ _00844_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10911__C1 _07250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout880 net881 vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08580__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15812_ net1197 vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__inv_2
Xfanout891 net895 vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12700__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16792_ clknet_leaf_38_wb_clk_i _02479_ _00775_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11824__B team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15743_ net1312 vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__inv_2
X_12955_ net1949 net870 net357 _03712_ vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_66_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11906_ net1754 net235 net479 vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__mux2_1
X_12886_ _05726_ net577 net360 vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__o21ba_1
XANTENNA__08883__A1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15674_ net1372 vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17413_ clknet_leaf_50_wb_clk_i _03100_ _01396_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_14625_ net1335 vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__inv_2
X_11837_ net2820 net243 net489 vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__mux2_1
XANTENNA__09013__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17344_ clknet_leaf_47_wb_clk_i _03031_ _01327_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_14556_ net1407 vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__inv_2
X_11768_ net2812 net201 net495 vssd1 vssd1 vccd1 vccd1 _03205_ sky130_fd_sc_hd__mux2_1
XANTENNA__09832__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17943__1458 vssd1 vssd1 vccd1 vccd1 _17943__1458/HI net1458 sky130_fd_sc_hd__conb_1
XANTENNA__09948__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14169__C1 net1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08852__C net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13507_ net185 _03964_ _03965_ net724 vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__a211o_1
X_10719_ _07001_ _07008_ net534 vssd1 vssd1 vccd1 vccd1 _07059_ sky130_fd_sc_hd__mux2_1
XANTENNA__12147__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14487_ net1399 vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__inv_2
X_17275_ clknet_leaf_69_wb_clk_i _02962_ _01258_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11699_ net1976 net284 net500 vssd1 vssd1 vccd1 vccd1 _03227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16226_ clknet_leaf_140_wb_clk_i net1642 _00214_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__dfrtp_1
X_13438_ _03889_ _03891_ _03897_ _03898_ _03885_ vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__o32a_1
XFILLER_0_130_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11986__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16157_ clknet_leaf_131_wb_clk_i _01920_ _00145_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13369_ net586 net565 team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1
+ vccd1 _03837_ sky130_fd_sc_hd__o21a_1
XANTENNA__11942__A1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15108_ net1233 vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__inv_2
X_16088_ clknet_leaf_132_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[10\]
+ _00076_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[10\] sky130_fd_sc_hd__dfrtp_1
X_15039_ net1314 vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09600_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[24\] net805 net777 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_127_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12610__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09531_ net1153 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[28\] net976
+ vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09462_ _05788_ _05791_ _05801_ net703 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__o32a_2
XFILLER_0_149_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08413_ net718 _04751_ vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__nor2_2
XFILLER_0_148_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09393_ _05570_ _05620_ _05658_ net559 vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__a31o_1
XFILLER_0_58_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout246_A _07842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08344_ net991 net948 vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__and2_1
XANTENNA__15222__A net1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12057__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08275_ net2352 net2109 net1042 vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout413_A _03563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1155_A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11896__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11749__X _07937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1322_A net1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout782_A net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12910__B1_N net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13135__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13964__X _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1108 net1114 vssd1 vssd1 vccd1 vccd1 net1108 sky130_fd_sc_hd__buf_1
XANTENNA__11146__C1 _07238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1119 net1120 vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_35_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09890__A net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09354__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout570_X net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout668_X net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11161__A2 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout187 _07639_ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_87_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12520__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout198 _07633_ vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09106__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08937__C net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09729_ _06066_ _06067_ net508 vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__a21boi_1
Xclkbuf_leaf_151_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_151_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13989__A2 _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout835_X net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12740_ net1598 net641 net609 _03587_ vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_83_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ net3021 net231 net389 vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ net1323 vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11622_ net3062 net216 net501 vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15390_ net1316 vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__inv_2
XANTENNA__09814__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10547__Y _06887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08672__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09130__A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14341_ net1338 vssd1 vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__inv_2
X_11553_ net1554 net1174 net590 vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10975__A2 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17060_ clknet_leaf_84_wb_clk_i _02747_ _01043_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10504_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[31\] net807 net755 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[31\]
+ _06832_ vssd1 vssd1 vccd1 vccd1 _06844_ sky130_fd_sc_hd__a221o_1
XFILLER_0_123_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14272_ net1340 vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__inv_2
X_11484_ net367 _07769_ net2052 net876 vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_107_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16011_ net1348 vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13223_ team_01_WB.instance_to_wrap.cpu.f0.num\[27\] net352 net348 net1906 vssd1
+ vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10435_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[27\] net804 _06752_
+ _06753_ _06754_ vssd1 vssd1 vccd1 vccd1 _06775_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_59_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13154_ net1618 net847 net839 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[22\] vssd1
+ vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10366_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[17\] net763 net622 vssd1
+ vssd1 vccd1 vccd1 _06706_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13126__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12105_ net2438 net235 net455 vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__mux2_1
X_17962_ net1477 vssd1 vssd1 vccd1 vccd1 la_data_out[4] sky130_fd_sc_hd__buf_2
X_13085_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[1\] net2244 net866 vssd1 vssd1
+ vccd1 vccd1 _02040_ sky130_fd_sc_hd__mux2_1
X_10297_ _04883_ net329 _04919_ vssd1 vssd1 vccd1 vccd1 _06637_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_148_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16913_ clknet_leaf_113_wb_clk_i _02600_ _00896_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_12036_ net2305 net241 net465 vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__mux2_1
XANTENNA__09008__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17893_ net1515 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
X_16844_ clknet_leaf_149_wb_clk_i _02531_ _00827_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12430__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10360__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16775_ clknet_leaf_105_wb_clk_i _02462_ _00758_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13987_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[64\] _04233_ _04263_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[120\]
+ _04278_ vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__a221o_1
X_15726_ net1297 vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_122_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10112__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12938_ _03694_ _03701_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[11\] net1038
+ vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_122_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12937__Y _03701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15657_ net1287 vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__inv_2
X_12869_ _06881_ net578 net361 vssd1 vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_34_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14608_ net1328 vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13601__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09805__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15588_ net1219 vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08582__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17327_ clknet_leaf_35_wb_clk_i _03014_ _01310_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14539_ net1426 vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08060_ _04522_ _04532_ _04536_ vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_70_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17258_ clknet_leaf_33_wb_clk_i _02945_ _01241_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_148_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16209_ clknet_leaf_123_wb_clk_i _01969_ _00197_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_144_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17189_ clknet_leaf_52_wb_clk_i _02876_ _01172_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10179__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12605__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11915__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09584__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13117__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08962_ _05043_ _05301_ vssd1 vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__or2_1
XANTENNA__09336__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08893_ net1107 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[2\] net943 vssd1
+ vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__and3_1
XANTENNA__11745__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12340__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10351__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12891__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08757__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout363_A _03580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14093__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14093__B2 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09514_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[29\] net800 net785 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__a22o_1
XANTENNA__10654__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09445_ net1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[29\] net943
+ vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout530_A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08773__B _05112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09376_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[26\] _04776_ net673 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[26\]
+ _05715_ vssd1 vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16523__CLK clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10406__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17986__1501 vssd1 vssd1 vccd1 vccd1 _17986__1501/HI net1501 sky130_fd_sc_hd__conb_1
X_08327_ net1137 net976 vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__and2_4
XFILLER_0_90_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13959__X _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1060_X net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout416_X net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09885__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14148__A2 _04226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08258_ net2591 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[15\] net1048 vssd1 vssd1
+ vccd1 vccd1 _03429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout997_A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12515__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08189_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[92\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[84\]
+ net1044 vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__mux2_1
X_10220_ _06550_ _06552_ _06556_ _06559_ vssd1 vssd1 vccd1 vccd1 _06560_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_37_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09575__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout785_X net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10543__B _06882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13108__A0 team_01_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10151_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[11\] net790 net739 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06491_ sky130_fd_sc_hd__a22o_1
XANTENNA__13659__A1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09327__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10082_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[7\] net738 _06412_ _06418_
+ _06419_ vssd1 vssd1 vccd1 vccd1 _06422_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13854__B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout952_X net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17942__1457 vssd1 vssd1 vccd1 vccd1 _17942__1457/HI net1457 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_7_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13910_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[9\] _04207_ vssd1 vssd1 vccd1
+ vccd1 _04208_ sky130_fd_sc_hd__or2_1
XANTENNA__12250__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14890_ net1283 vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__inv_2
XANTENNA__12882__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08667__C net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13841_ net1179 net1066 net3180 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[2\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_69_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13772_ _04156_ _01836_ vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__or2_1
X_16560_ clknet_leaf_159_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[26\]
+ _00543_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10984_ _07277_ _07283_ net524 vssd1 vssd1 vccd1 vccd1 _07324_ sky130_fd_sc_hd__mux2_1
XANTENNA__08964__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10645__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15511_ net1243 vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__inv_2
X_12723_ net1032 team_01_WB.instance_to_wrap.cpu.f0.write_i vssd1 vssd1 vccd1 vccd1
+ _03574_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_100_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16491_ clknet_leaf_156_wb_clk_i _02245_ _00474_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_15442_ net1290 vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__inv_2
X_12654_ _07791_ _07793_ net573 vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__and3_4
X_11605_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[31\] _07821_ vssd1 vssd1
+ vccd1 vccd1 _07822_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12585_ net3076 net318 net402 vssd1 vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__mux2_1
X_15373_ net1267 vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17112_ clknet_leaf_49_wb_clk_i _02799_ _01095_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11536_ net1983 net1174 net589 net1163 vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__a22o_1
X_14324_ net1348 vssd1 vssd1 vccd1 vccd1 _00118_ sky130_fd_sc_hd__inv_2
XANTENNA__14139__A2 _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_59 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14255_ net1226 vssd1 vssd1 vccd1 vccd1 _00049_ sky130_fd_sc_hd__inv_2
X_17043_ clknet_leaf_17_wb_clk_i _02730_ _01026_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11467_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[29\] net579 vssd1 vssd1 vccd1
+ vccd1 _07761_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12425__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10734__A _06912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13206_ net33 net836 net629 net2077 vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10418_ net1132 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[27\] net948
+ vssd1 vssd1 vccd1 vccd1 _06758_ sky130_fd_sc_hd__and3b_1
X_14186_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[12\] _04453_ net1837 vssd1
+ vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__a21oi_1
X_11398_ _04468_ _07721_ _07722_ vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_74_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13137_ net1653 net846 net633 team_01_WB.instance_to_wrap.a1.ADR_I\[6\] vssd1 vssd1
+ vccd1 vccd1 _02004_ sky130_fd_sc_hd__a22o_1
X_10349_ net991 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[17\] net973 vssd1
+ vssd1 vccd1 vccd1 _06689_ sky130_fd_sc_hd__and3_1
XFILLER_0_104_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_146_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17945_ net1460 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
X_13068_ net2307 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[26\] net864 vssd1 vssd1
+ vccd1 vccd1 _02057_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12019_ net1829 net294 net468 vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__mux2_1
XANTENNA__12160__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_79_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17876_ clknet_leaf_131_wb_clk_i _03551_ _01816_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12873__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09035__A _05338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16827_ clknet_leaf_74_wb_clk_i _02514_ _00810_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10884__A1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10884__B2 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16758_ clknet_leaf_25_wb_clk_i _02445_ _00741_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10636__A1 _06919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15709_ net1313 vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__inv_2
X_16689_ clknet_leaf_116_wb_clk_i _02376_ _00672_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_146_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09230_ net376 _05378_ _05493_ _05569_ vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__and4_1
XFILLER_0_150_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11079__A_N net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_14_Left_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09161_ net1091 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[16\] net927
+ vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__and3_1
XANTENNA__09254__A1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09201__C net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10347__C net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08112_ _04480_ team_01_WB.instance_to_wrap.cpu.f0.num\[14\] team_01_WB.instance_to_wrap.cpu.f0.num\[9\]
+ _04484_ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__a22o_1
X_09092_ net1012 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[13\] net882 vssd1
+ vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17695__Q team_01_WB.instance_to_wrap.cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_141_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08043_ net1661 net570 net347 team_01_WB.instance_to_wrap.cpu.f0.i\[12\] vssd1 vssd1
+ vccd1 vccd1 _03548_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold900 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2435 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12335__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold911 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2446 sky130_fd_sc_hd__dlygate4sd3_1
Xhold922 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[97\] vssd1 vssd1 vccd1 vccd1
+ net2457 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout209_A _07847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09557__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold933 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2468 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08114__A team_01_WB.instance_to_wrap.cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_40_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold944 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold955 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[67\] vssd1 vssd1 vccd1 vccd1
+ net2490 sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2501 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16104__Q team_01_WB.instance_to_wrap.cpu.f0.data_adr\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold977 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2512 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_23_Left_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09994_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[2\] _04636_ net813 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06334_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1020_A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold988 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2523 sky130_fd_sc_hd__dlygate4sd3_1
Xhold999 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2534 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09309__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08945_ net1027 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[6\] net903 vssd1
+ vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_32_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout480_A _07949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1600 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net3135 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1611 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net3146 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12070__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08876_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[3\] _04771_ _05199_ _05203_
+ _05205_ vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__a2111o_1
Xhold1622 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 net3157
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1633 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net3168 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09319__A_N _04844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1644 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 net3179
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout745_A net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout912_A net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout533_X net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10819__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09428_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[28\] net662 net648 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05768_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout700_X net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09359_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[25\] net689 _04778_
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[25\] vssd1 vssd1 vccd1 vccd1
+ _05699_ sky130_fd_sc_hd__a22o_1
XANTENNA__08048__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09796__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12370_ net2957 net237 net423 vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11321_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[6\] net1176 _04534_ _07652_ vssd1
+ vssd1 vccd1 vccd1 _07657_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12245__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14040_ net147 net604 vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_95_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11252_ _05681_ _06919_ net511 vssd1 vssd1 vccd1 vccd1 _07592_ sky130_fd_sc_hd__or3b_1
X_10203_ net1140 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[8\] _04662_
+ vssd1 vssd1 vccd1 vccd1 _06543_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_113_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11183_ net337 _07376_ _07522_ vssd1 vssd1 vccd1 vccd1 _07523_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_52_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input41_A wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10134_ net1144 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[11\] net972
+ vssd1 vssd1 vccd1 vccd1 _06474_ sky130_fd_sc_hd__and3_1
X_15991_ net1413 vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__inv_2
X_17730_ clknet_leaf_123_wb_clk_i _03406_ _01670_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10065_ _06313_ _06315_ vssd1 vssd1 vccd1 vccd1 _06405_ sky130_fd_sc_hd__xor2_2
X_14942_ net1316 vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_141_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17906__1441 vssd1 vssd1 vccd1 vccd1 _17906__1441/HI net1441 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_141_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10866__A1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17661_ clknet_leaf_3_wb_clk_i _03346_ _01602_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09720__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14873_ net1231 vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__inv_2
XANTENNA__14057__A1 team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16612_ clknet_leaf_82_wb_clk_i _02299_ _00595_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13824_ net3073 net832 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[17\]
+ sky130_fd_sc_hd__and2_1
X_17592_ clknet_leaf_89_wb_clk_i _03279_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16543_ clknet_leaf_6_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[9\]
+ _00526_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13755_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[7\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[6\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__or4b_1
X_10967_ net343 _07294_ _07305_ _07071_ vssd1 vssd1 vccd1 vccd1 _07307_ sky130_fd_sc_hd__o22a_1
XANTENNA__10729__A _06920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12706_ net1911 net255 net384 vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__mux2_1
XANTENNA__10094__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11291__A1 _06886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16474_ clknet_leaf_140_wb_clk_i _02228_ _00457_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10898_ net530 _07237_ _07235_ vssd1 vssd1 vccd1 vccd1 _07238_ sky130_fd_sc_hd__a21boi_2
X_13686_ team_01_WB.instance_to_wrap.cpu.c0.count\[14\] team_01_WB.instance_to_wrap.cpu.c0.count\[13\]
+ _04108_ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15425_ net1281 vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__inv_2
XANTENNA__09021__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12637_ net2040 net263 net393 vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13742__A_N net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_152_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12568_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[19\] net239 net399 vssd1
+ vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__mux2_1
X_15356_ net1249 vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_117_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09956__C net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08860__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_152_Right_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14307_ net1324 vssd1 vssd1 vccd1 vccd1 _00101_ sky130_fd_sc_hd__inv_2
XANTENNA__13111__Y _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11519_ team_01_WB.instance_to_wrap.cpu.DM0.enable net714 vssd1 vssd1 vccd1 vccd1
+ _07783_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12155__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12499_ net2081 net201 net407 vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15287_ net1215 vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold207 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[122\] vssd1 vssd1 vccd1 vccd1
+ net1742 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold218 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1753 sky130_fd_sc_hd__dlygate4sd3_1
X_17026_ clknet_leaf_75_wb_clk_i _02713_ _01009_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold229 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[12\] vssd1 vssd1 vccd1 vccd1 net1764
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14238_ net1336 vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__inv_2
XANTENNA__12950__Y _03710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11994__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14169_ net1823 _04189_ _04445_ net1426 vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_21_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09317__X _05657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11295__A net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08730_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[5\] net676 _05060_ net706
+ vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__a211o_1
X_17928_ net1535 vssd1 vssd1 vccd1 vccd1 gpio_oeb[37] sky130_fd_sc_hd__buf_2
X_17985__1500 vssd1 vssd1 vccd1 vccd1 _17985__1500/HI net1500 sky130_fd_sc_hd__conb_1
XFILLER_0_56_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1280 net1281 vssd1 vssd1 vccd1 vccd1 net1280 sky130_fd_sc_hd__buf_4
Xfanout1291 net1292 vssd1 vssd1 vccd1 vccd1 net1291 sky130_fd_sc_hd__buf_4
X_08661_ _04997_ _04998_ _04999_ _05000_ vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__or4_2
XANTENNA__10857__A1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09711__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17859_ clknet_leaf_138_wb_clk_i _03534_ _01799_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.read_i
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10857__B2 _04970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08592_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[15\] net685 net662 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__a22o_1
XANTENNA__10609__A1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10085__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08109__A _04504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09213_ net1085 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[17\] net882
+ vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__and3_1
XFILLER_0_147_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10077__C net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17941__1456 vssd1 vssd1 vccd1 vccd1 _17941__1456/HI net1456 sky130_fd_sc_hd__conb_1
X_09144_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[14\] net682 _05464_
+ _05466_ _05471_ vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_20_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09075_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[12\] net704 _05411_ _05414_
+ vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_32_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12065__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1235_A net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08026_ team_01_WB.instance_to_wrap.cpu.K0.code\[2\] _04521_ team_01_WB.instance_to_wrap.cpu.K0.code\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__or3b_2
XFILLER_0_102_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold730 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2265 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold741 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[31\] vssd1 vssd1 vccd1 vccd1
+ net2276 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold752 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2287 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold763 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold774 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2320 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1402_A net1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold796 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2331 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09977_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[2\] net798 _04659_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06317_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout483_X net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout862_A net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13972__X _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08928_ net1027 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[6\] net915 vssd1
+ vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__and3_1
XFILLER_0_99_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1430 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2965 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1441 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2976 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10848__A1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1452 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[6\] vssd1 vssd1 vccd1 vccd1
+ net2987 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout650_X net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08859_ net1024 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[3\] net915 vssd1
+ vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__and3_1
Xhold1463 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2998 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12588__X _03567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout748_X net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1474 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net3009 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1485 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[104\] vssd1 vssd1 vccd1 vccd1
+ net3020 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1496 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net3031 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_58_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11870_ net2253 net241 net485 vssd1 vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__mux2_1
XANTENNA__08945__C net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10821_ net528 _07068_ _07159_ vssd1 vssd1 vccd1 vccd1 _07161_ sky130_fd_sc_hd__a21o_1
XANTENNA__11652__B net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout915_X net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10752_ _06001_ _06034_ _07091_ vssd1 vssd1 vccd1 vccd1 _07092_ sky130_fd_sc_hd__or3_1
X_13540_ _03926_ _03992_ vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__xor2_1
XFILLER_0_137_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13471_ _03930_ _03931_ vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__and2_1
X_10683_ net537 _07022_ net548 vssd1 vssd1 vccd1 vccd1 _07023_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_97_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12422_ net2273 net289 net420 vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__mux2_1
X_15210_ net1385 vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_97_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09769__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16190_ clknet_leaf_1_wb_clk_i _01950_ _00178_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08306__X _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08680__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12773__A1 _07251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15141_ net1262 vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__inv_2
X_12353_ net2002 net305 net430 vssd1 vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11304_ _07642_ _07643_ vssd1 vssd1 vccd1 vccd1 _07644_ sky130_fd_sc_hd__xnor2_1
X_15072_ net1272 vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__inv_2
X_12284_ net3167 net299 net438 vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12525__A1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14023_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[34\] _04221_ _04233_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[66\]
+ vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__a22o_1
X_11235_ net369 _07348_ _07349_ net336 _07574_ vssd1 vssd1 vccd1 vccd1 _07575_ sky130_fd_sc_hd__a221o_1
XFILLER_0_121_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12703__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10536__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08689__A net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11166_ net558 _07499_ _07505_ _07071_ vssd1 vssd1 vccd1 vccd1 _07506_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_101_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10117_ _06445_ _06448_ _06453_ _06456_ vssd1 vssd1 vccd1 vccd1 _06457_ sky130_fd_sc_hd__or4_1
XFILLER_0_140_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15974_ net1405 vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__inv_2
X_11097_ _06901_ _06913_ _07436_ vssd1 vssd1 vccd1 vccd1 _07437_ sky130_fd_sc_hd__or3_1
XANTENNA__10450__C net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17713_ clknet_leaf_125_wb_clk_i _03397_ _01654_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14925_ net1264 vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__inv_2
X_10048_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[0\] net807 net772 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06388_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_3_4_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09016__C net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold90 team_01_WB.instance_to_wrap.cpu.f0.write_data\[30\] vssd1 vssd1 vccd1 vccd1
+ net1625 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11500__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17644_ clknet_leaf_157_wb_clk_i _03329_ _01585_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.bit30
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_69_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14856_ net1375 vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__inv_2
XANTENNA__08855__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13807_ net1711 net832 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[0\]
+ sky130_fd_sc_hd__and2_1
X_17575_ clknet_leaf_122_wb_clk_i _03262_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__dfxtp_1
X_14787_ net1218 vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11999_ net2889 net208 net468 vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16526_ clknet_leaf_0_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[24\]
+ _00509_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13738_ team_01_WB.instance_to_wrap.cpu.DM0.dhit net1176 vssd1 vssd1 vccd1 vccd1
+ team_01_WB.instance_to_wrap.cpu.f0.next_lcd_en sky130_fd_sc_hd__and2_1
XFILLER_0_46_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11989__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16457_ clknet_leaf_16_wb_clk_i _02211_ _00440_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13669_ net1178 _03735_ _04099_ vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15408_ net1279 vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16388_ clknet_leaf_96_wb_clk_i net2338 _00371_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[111\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12764__A1 _07621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15339_ net1425 vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09900_ _06236_ _06237_ _06238_ _06239_ vssd1 vssd1 vccd1 vccd1 _06240_ sky130_fd_sc_hd__or4_1
X_17009_ clknet_leaf_115_wb_clk_i _02696_ _00992_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12613__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10527__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09393__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09831_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[13\] net791 net733 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06171_ sky130_fd_sc_hd__a22o_1
Xfanout517 net518 vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout528 net529 vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__clkbuf_4
Xfanout539 net541 vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__clkbuf_4
X_09762_ _06002_ _06036_ _06068_ _06101_ vssd1 vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__or4_1
X_08713_ net1097 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[5\] net898 vssd1
+ vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__and3_1
X_09693_ _05657_ _05732_ vssd1 vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__xnor2_1
X_08644_ net1102 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[10\] net898
+ vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08575_ net1000 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[19\] net940 vssd1
+ vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__and3_1
XANTENNA__10369__A _04970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout443_A _07959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10058__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09999__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08120__B2 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11899__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1352_A net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13399__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09596__C net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09127_ net1109 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[14\] net916
+ vssd1 vssd1 vccd1 vccd1 _05467_ sky130_fd_sc_hd__and3_1
XANTENNA__13967__X _04259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17905__1440 vssd1 vssd1 vccd1 vccd1 _17905__1440/HI net1440 sky130_fd_sc_hd__conb_1
XANTENNA__12871__X _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_105_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_105_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_92_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09058_ net1113 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[12\] net941
+ vssd1 vssd1 vccd1 vccd1 _05398_ sky130_fd_sc_hd__and3_1
XANTENNA__09893__A net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout698_X net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08009_ team_01_WB.instance_to_wrap.cpu.K0.keyvalid vssd1 vssd1 vccd1 vccd1 _04506_
+ sky130_fd_sc_hd__inv_2
Xhold560 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2095 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12523__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold571 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[14\] vssd1 vssd1 vccd1 vccd1
+ net2106 sky130_fd_sc_hd__dlygate4sd3_1
Xhold582 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2117 sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ _05529_ net371 vssd1 vssd1 vccd1 vccd1 _07360_ sky130_fd_sc_hd__nor2_1
Xhold593 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2128 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08302__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_10__f_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11366__C net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08021__B _04516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10270__C net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12971_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[115\] net1788 net861 vssd1 vssd1
+ vccd1 vccd1 _02154_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1260 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2795 sky130_fd_sc_hd__dlygate4sd3_1
X_14710_ net1193 vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__inv_2
Xhold1271 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2806 sky130_fd_sc_hd__dlygate4sd3_1
X_11922_ net2164 net320 net482 vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__mux2_1
Xhold1282 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2817 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1293 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[55\] vssd1 vssd1 vccd1 vccd1
+ net2828 sky130_fd_sc_hd__dlygate4sd3_1
X_15690_ net1283 vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08675__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09133__A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14641_ net1378 vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11853_ net1897 net292 net490 vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__mux2_1
XANTENNA__10049__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10804_ _06919_ _07143_ vssd1 vssd1 vccd1 vccd1 _07144_ sky130_fd_sc_hd__nor2_1
XANTENNA__11246__A1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17360_ clknet_leaf_145_wb_clk_i _03047_ _01343_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_11784_ net2209 net298 net497 vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14572_ net1421 vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16311_ clknet_leaf_102_wb_clk_i _02065_ _00294_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13523_ net187 _03977_ _03978_ net727 vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_136_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10735_ _05781_ net331 _07073_ net334 net370 vssd1 vssd1 vccd1 vccd1 _07075_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17291_ clknet_leaf_9_wb_clk_i _02978_ _01274_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09787__B net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08662__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16242_ clknet_leaf_151_wb_clk_i net1570 _00230_ vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__dfrtp_1
X_13454_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] _05495_ vssd1 vssd1
+ vccd1 vccd1 _03915_ sky130_fd_sc_hd__or2_1
X_10666_ net551 _06313_ _07005_ vssd1 vssd1 vccd1 vccd1 _07006_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12405_ net2126 net268 net420 vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13385_ _03845_ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__inv_2
X_16173_ clknet_leaf_6_wb_clk_i _01933_ _00161_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10597_ net374 _06158_ net544 vssd1 vssd1 vccd1 vccd1 _06937_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10445__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15124_ net1378 vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__inv_2
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__buf_2
X_12336_ net3011 net269 net427 vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12941__B net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15055_ net1388 vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__inv_2
XANTENNA__12433__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12267_ net2263 net205 net435 vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14006_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[81\] _04251_ _04260_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[57\]
+ _04296_ vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__a221o_1
X_11218_ net504 net333 net331 vssd1 vssd1 vccd1 vccd1 _07558_ sky130_fd_sc_hd__a21o_1
XANTENNA__09375__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12198_ net1989 net273 net445 vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__mux2_1
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__buf_2
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__buf_2
XFILLER_0_128_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11721__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11149_ _07482_ _07486_ _07488_ vssd1 vssd1 vccd1 vccd1 _07489_ sky130_fd_sc_hd__or3_4
XANTENNA__14120__B1 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13930__A_N team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15957_ net1418 vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_108_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17940__1455 vssd1 vssd1 vccd1 vccd1 _17940__1455/HI net1455 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_108_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10288__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14908_ net1244 vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__inv_2
X_15888_ net1399 vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__inv_2
XANTENNA__08585__C net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17627_ clknet_leaf_3_wb_clk_i _03312_ _01568_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_59_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14839_ net1243 vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__inv_2
XANTENNA__09978__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08360_ _04696_ _04697_ _04698_ _04699_ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__or4_1
X_17558_ clknet_leaf_29_wb_clk_i _03245_ _01541_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_3_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16509_ clknet_leaf_6_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[7\]
+ _00492_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_08291_ net1158 net1164 net1166 net1161 vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_156_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12608__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17489_ clknet_leaf_143_wb_clk_i _03176_ _01472_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09850__A1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10996__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11512__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09189__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10460__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_6__f_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10212__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12343__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout303 _07912_ vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09905__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout314 net315 vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__clkbuf_2
Xfanout325 net326 vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__buf_1
XANTENNA_fanout393_A net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16112__Q team_01_WB.instance_to_wrap.cpu.f0.data_adr\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout336 net337 vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__buf_2
X_09814_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[14\] net809 net792 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06154_ sky130_fd_sc_hd__a22o_1
Xfanout347 _04526_ vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__buf_4
Xfanout358 net359 vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09381__A3 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1100_A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout369 net370 vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14111__B1 _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09745_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[20\] net739 _06071_ _06077_
+ _06081_ vssd1 vssd1 vccd1 vccd1 _06085_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_20_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout560_A net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout658_A _04813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08877__C1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09676_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[22\] net776 net734 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06016_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_6_Left_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08627_ _04952_ _04963_ _04964_ _04966_ vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__or4_1
XFILLER_0_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout446_X net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout825_A _04579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1090_X net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09888__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08558_ net999 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[19\] net925 vssd1
+ vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__and3_1
XFILLER_0_83_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12518__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08489_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[23\] net690 _04777_ _04792_
+ _04764_ vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_37_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1355_X net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10520_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[31\] net687 net684 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06860_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10451_ net1147 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[26\] net952
+ vssd1 vssd1 vccd1 vccd1 _06791_ sky130_fd_sc_hd__and3b_1
XFILLER_0_91_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10265__C net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13170_ net1922 net848 net840 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[6\] vssd1
+ vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10382_ net994 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[16\] net945 vssd1
+ vssd1 vccd1 vccd1 _06722_ sky130_fd_sc_hd__o21a_1
XANTENNA__13857__B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout982_X net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12121_ net2830 net318 net458 vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12253__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09357__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12052_ net2764 net293 net466 vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__mux2_1
Xhold390 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1925 sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ _05758_ net504 vssd1 vssd1 vccd1 vccd1 _07343_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_73_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16860_ clknet_leaf_60_wb_clk_i _02547_ _00843_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10911__B1 _07239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout870 net871 vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__clkbuf_4
X_15811_ net1197 vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__inv_2
XANTENNA__14102__B1 _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout881 _04810_ vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__clkbuf_4
Xfanout892 net895 vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__clkbuf_4
X_16791_ clknet_leaf_13_wb_clk_i _02478_ _00774_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_29_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15742_ net1318 vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__inv_2
X_12954_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[5\] _05074_ net1038 vssd1
+ vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2625 sky130_fd_sc_hd__dlygate4sd3_1
X_11905_ net1967 net239 net479 vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__mux2_1
X_15673_ net1232 vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__inv_2
XANTENNA_output110_A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12885_ net1846 net872 net359 _03664_ vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__a22o_1
XANTENNA__08883__A2 _05219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17412_ clknet_leaf_82_wb_clk_i _03099_ _01395_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ net1337 vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__inv_2
X_11836_ net2210 net201 net487 vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_155_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ clknet_leaf_44_wb_clk_i _03030_ _01326_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14555_ net1427 vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__inv_2
XANTENNA__10296__X _06636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10978__A0 _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12428__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11767_ net2243 net203 net495 vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__mux2_1
X_13506_ net198 net194 _07830_ net644 vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17274_ clknet_leaf_76_wb_clk_i _02961_ _01257_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10718_ _06998_ _07002_ net534 vssd1 vssd1 vccd1 vccd1 _07058_ sky130_fd_sc_hd__mux2_1
X_14486_ net1351 vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11698_ net614 _07807_ _07895_ _07894_ vssd1 vssd1 vccd1 vccd1 _07896_ sky130_fd_sc_hd__a31o_4
XFILLER_0_55_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16225_ clknet_leaf_140_wb_clk_i net1612 _00213_ vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__dfrtp_1
X_13437_ team_01_WB.instance_to_wrap.cpu.CU0.bit30 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\]
+ net595 _03886_ vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10649_ net511 net510 net543 vssd1 vssd1 vccd1 vccd1 _06989_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08399__A1 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16156_ clknet_leaf_134_wb_clk_i _01919_ _00144_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13368_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[9\] _04579_ _07650_ _03836_
+ vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__o22a_1
X_15107_ net1220 vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__inv_2
X_12319_ net2023 net310 net431 vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__mux2_1
XANTENNA__12163__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16087_ clknet_leaf_132_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[9\]
+ _00075_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[9\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10472__A _06811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13299_ _04516_ _03745_ _03782_ team_01_WB.instance_to_wrap.cpu.f0.next_write_i vssd1
+ vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__o31a_1
XANTENNA__09348__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15038_ net1316 vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_127_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16989_ clknet_leaf_75_wb_clk_i _02676_ _00972_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09530_ net513 _05868_ vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09461_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[29\] net653 _05795_
+ _05799_ _05800_ vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09204__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08874__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08412_ _04708_ net725 net718 vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__or3_4
X_09392_ _05570_ _05620_ net559 vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12958__A1 _05219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08343_ net995 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[30\] net963 vssd1
+ vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12338__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08626__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08274_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[7\] net1537 net1042 vssd1 vssd1
+ vccd1 vccd1 _03413_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08117__A team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_104_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout406_A _03565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1148_A net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11394__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_70_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12073__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1315_A net1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1109 net1114 vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout396_X net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout775_A _04667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12801__S net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1103_X net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08787__A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout188 net191 vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_87_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout942_A _04759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout199 _07633_ vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_87_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07989_ team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1 _04487_
+ sky130_fd_sc_hd__inv_2
XANTENNA_fanout563_X net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11449__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09728_ net508 _06066_ _06067_ vssd1 vssd1 vccd1 vccd1 _06068_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_83_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout730_X net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09659_ net510 _05998_ vssd1 vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__nand2_1
X_12670_ net2091 net262 net388 vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11621_ _07832_ _07834_ net612 vssd1 vssd1 vccd1 vccd1 _07835_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_13_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12248__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_120_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_120_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10557__A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08617__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14340_ net1338 vssd1 vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__inv_2
XANTENNA__10424__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11552_ net1553 net1173 net590 vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10975__A3 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10503_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[31\] net817 net779 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06843_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_150_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11483_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[21\] net580 vssd1 vssd1 vccd1
+ vccd1 _07769_ sky130_fd_sc_hd__nand2_1
X_14271_ net1342 vssd1 vssd1 vccd1 vccd1 _00065_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16010_ net1357 vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13222_ team_01_WB.instance_to_wrap.cpu.f0.num\[28\] net352 net348 team_01_WB.instance_to_wrap.cpu.f0.i\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__a22o_1
XANTENNA_input71_A wbs_cyc_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10434_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[27\] net777 net730 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06774_ sky130_fd_sc_hd__a22o_1
XANTENNA__13374__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_150_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08314__X _04654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10563__Y _06903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13079__S net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10365_ net769 _06697_ _06701_ _06704_ vssd1 vssd1 vccd1 vccd1 _06705_ sky130_fd_sc_hd__nor4_1
X_13153_ net1603 net847 net839 net1587 vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_5__f_wb_clk_i_X clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12104_ net3063 net237 net455 vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__mux2_1
X_17961_ net1476 vssd1 vssd1 vccd1 vccd1 la_data_out[3] sky130_fd_sc_hd__buf_2
X_13084_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[2\] net2398 net864 vssd1 vssd1
+ vccd1 vccd1 _02041_ sky130_fd_sc_hd__mux2_1
X_10296_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] net625 _06634_ _06635_
+ vssd1 vssd1 vccd1 vccd1 _06636_ sky130_fd_sc_hd__a22o_2
XANTENNA__11137__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08538__D1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12035_ net2345 _07858_ net464 vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__mux2_1
XANTENNA__11328__A_N team_01_WB.instance_to_wrap.cpu.DM0.data_i\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16912_ clknet_leaf_146_wb_clk_i _02599_ _00895_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11688__A1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12711__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17892_ net1514 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
XANTENNA__12885__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_69_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09750__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16843_ clknet_leaf_8_wb_clk_i _02530_ _00826_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_69_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16774_ clknet_leaf_74_wb_clk_i _02461_ _00757_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13986_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[8\] _04253_ _04264_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[104\]
+ vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__a22o_1
X_15725_ net1264 vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__inv_2
X_12937_ _04968_ _07756_ vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_122_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08856__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15656_ net1375 vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__inv_2
X_12868_ _04753_ _04944_ _07630_ net578 _03652_ vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__o311a_1
XFILLER_0_68_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08863__C net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14607_ net1328 vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11819_ net2411 net310 net491 vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__mux2_1
XANTENNA__12158__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15587_ net1221 vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__inv_2
X_12799_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] net1060 net362 _03627_
+ vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17326_ clknet_leaf_27_wb_clk_i _03013_ _01309_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14538_ net1366 vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_78_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11997__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17257_ clknet_leaf_39_wb_clk_i _02944_ _01240_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_895 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14469_ net1356 vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__inv_2
X_16208_ clknet_leaf_123_wb_clk_i _01968_ _00196_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__dfrtp_1
X_17188_ clknet_leaf_73_wb_clk_i _02875_ _01171_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09033__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16139_ clknet_leaf_131_wb_clk_i _01902_ _00127_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08961_ net602 _05300_ _05266_ vssd1 vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__a21o_2
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08892_ net1025 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[2\] net941 vssd1
+ vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__and3_1
XANTENNA__12876__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Left_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11745__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08400__A team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14093__A2 _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09513_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[29\] net757 net735 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10929__X _07269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11300__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout356_A _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1098_A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09444_ net1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[29\] net881
+ vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13589__D1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09231__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10377__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09375_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[26\] _04778_ net677 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__a22o_1
XANTENNA__12068__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_96_Left_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08326_ net1155 net949 vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09272__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08257_ net2816 net2572 net1046 vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout409_X net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08188_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[93\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[85\]
+ net1050 vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__mux2_1
XANTENNA__09024__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout892_A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10824__B net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13975__X _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_103_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13108__A1 net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09980__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10150_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[11\] net794 _06487_ _06488_
+ _06489_ vssd1 vssd1 vccd1 vccd1 _06490_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout680_X net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout778_X net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10081_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[7\] net799 net736 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06421_ sky130_fd_sc_hd__a22o_1
XANTENNA__12531__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08948__C net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout945_X net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13840_ net1179 net1066 net3173 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[1\]
+ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_18_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14084__A2 _04221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13771_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[3\] _04152_ _04157_ net1183
+ vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__o211a_1
X_10983_ _07316_ _07322_ _07310_ vssd1 vssd1 vccd1 vccd1 _07323_ sky130_fd_sc_hd__or3b_4
X_15510_ net1256 vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12722_ net1170 _04718_ team_01_WB.instance_to_wrap.cpu.DM0.enable team_01_WB.instance_to_wrap.cpu.DM0.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__or4b_1
X_16490_ clknet_leaf_152_wb_clk_i _02244_ _00473_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08309__X _04649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08683__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_133_Right_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15441_ net1420 vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__inv_2
X_12653_ net2070 net289 net394 vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09799__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11604_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\]
+ _07820_ vssd1 vssd1 vccd1 vccd1 _07821_ sky130_fd_sc_hd__and3_1
XANTENNA__13595__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15372_ net1260 vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__inv_2
X_12584_ net2424 net305 net401 vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_142_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_25_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09263__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17111_ clknet_leaf_16_wb_clk_i _02798_ _01094_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14323_ net1329 vssd1 vssd1 vccd1 vccd1 _00117_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11535_ net2627 net1172 net589 net1160 vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__a22o_1
XANTENNA__11070__A2 _06526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12706__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17042_ clknet_leaf_143_wb_clk_i _02729_ _01025_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input74_X net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14254_ net1226 vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_78_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11466_ net366 _07760_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[30\] net874
+ vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_78_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13205_ net3 net837 _03738_ net3075 vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__a22o_1
X_10417_ net1132 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[27\] net956
+ vssd1 vssd1 vccd1 vccd1 _06757_ sky130_fd_sc_hd__and3_1
X_14185_ net2903 _04453_ _04455_ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__o21a_1
X_11397_ _07668_ _07696_ _07714_ net1068 vssd1 vssd1 vccd1 vccd1 _07722_ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10453__C net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08774__A1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13136_ net1622 net845 net633 team_01_WB.instance_to_wrap.a1.ADR_I\[7\] vssd1 vssd1
+ vccd1 vccd1 _02005_ sky130_fd_sc_hd__a22o_1
X_10348_ net1139 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[17\] net980
+ vssd1 vssd1 vccd1 vccd1 _06688_ sky130_fd_sc_hd__and3_1
XFILLER_0_104_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09019__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15318__A net1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12441__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17944_ net1459 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
X_10279_ net1128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[19\] net972
+ vssd1 vssd1 vccd1 vccd1 _06619_ sky130_fd_sc_hd__and3_1
X_13067_ net3015 net2958 net861 vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__mux2_1
X_12018_ net2822 net298 net469 vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__mux2_1
XANTENNA__08858__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17875_ clknet_leaf_138_wb_clk_i _03550_ _01815_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_46 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16826_ clknet_leaf_80_wb_clk_i _02513_ _00809_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11284__C _07621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14075__A2 _04246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16757_ clknet_leaf_111_wb_clk_i _02444_ _00740_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13969_ _04218_ _04224_ vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__nor2_4
XANTENNA__11581__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15708_ net1245 vssd1 vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__inv_2
XANTENNA__11294__C1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16688_ clknet_leaf_146_wb_clk_i _02375_ _00671_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15639_ net1214 vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09160_ net1010 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[16\] net940 vssd1
+ vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__and3_1
XFILLER_0_57_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09254__A2 _05591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08111_ net1070 team_01_WB.instance_to_wrap.cpu.f0.num\[8\] vssd1 vssd1 vccd1 vccd1
+ _04581_ sky130_fd_sc_hd__and2_1
XFILLER_0_145_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17309_ clknet_leaf_69_wb_clk_i _02996_ _01292_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09091_ net1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[13\] net944
+ vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12616__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08042_ net1600 net570 net346 team_01_WB.instance_to_wrap.cpu.f0.i\[13\] vssd1 vssd1
+ vccd1 vccd1 _03549_ sky130_fd_sc_hd__a22o_1
XANTENNA__11299__Y _07639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold901 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2436 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold912 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2447 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold923 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2458 sky130_fd_sc_hd__dlygate4sd3_1
Xhold934 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2469 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09411__C1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold945 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[51\] vssd1 vssd1 vccd1 vccd1
+ net2480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold956 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2491 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10021__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09962__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold967 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2502 sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2513 sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ _06320_ _06324_ _06329_ _06332_ vssd1 vssd1 vccd1 vccd1 _06333_ sky130_fd_sc_hd__or4_1
Xhold989 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2524 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15228__A net1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08944_ net1111 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[6\] net931 vssd1
+ vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__and3_1
XANTENNA__12351__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1013_A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1601 team_01_WB.instance_to_wrap.cpu.f0.num\[6\] vssd1 vssd1 vccd1 vccd1 net3136
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09714__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1612 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net3147 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08875_ _05209_ _05210_ _05213_ _05214_ vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_4_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1623 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[13\] vssd1 vssd1 vccd1 vccd1 net3158
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout473_A _07952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1634 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net3169 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09190__A1 net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16120__Q team_01_WB.instance_to_wrap.cpu.f0.data_adr\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold1645 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 net3180
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout640_A _03572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1382_A net1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout359_X net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09599__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08150__C1 _04516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09493__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09427_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[28\] net695 net676 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[28\]
+ _05766_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout905_A net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13577__A1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09358_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[25\] net665 net706 vssd1
+ vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08309_ net1139 net968 vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__and2_4
XFILLER_0_74_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09289_ net1004 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[22\] net923 vssd1
+ vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__and3_1
XANTENNA__12526__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11320_ _07656_ net1537 _07655_ vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout895_X net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11251_ net336 _07351_ vssd1 vssd1 vccd1 vccd1 _07591_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_95_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10273__C net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10012__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10202_ net992 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[8\] net968 vssd1
+ vssd1 vccd1 vccd1 _06542_ sky130_fd_sc_hd__and3_1
XANTENNA__09953__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11182_ _05006_ net330 _07376_ _06919_ _06915_ vssd1 vssd1 vccd1 vccd1 _07522_ sky130_fd_sc_hd__o221a_1
X_10133_ net1144 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[11\] net956
+ vssd1 vssd1 vccd1 vccd1 _06473_ sky130_fd_sc_hd__and3_1
XANTENNA__12261__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15990_ net1407 vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__inv_2
XANTENNA__08678__C net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13501__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input34_A gpio_in[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ _06402_ _06403_ _06343_ vssd1 vssd1 vccd1 vccd1 _06404_ sky130_fd_sc_hd__a21o_1
X_14941_ net1236 vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_141_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17660_ clknet_leaf_3_wb_clk_i _03345_ _01601_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_141_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14872_ net1209 vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16611_ clknet_leaf_63_wb_clk_i _02298_ _00594_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13823_ net1655 net832 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[16\]
+ sky130_fd_sc_hd__and2_1
X_17591_ clknet_leaf_129_wb_clk_i _03278_ _01550_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.code\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13092__S net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16542_ clknet_leaf_5_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[8\]
+ _00525_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13754_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[8\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[13\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[12\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__or4b_1
XFILLER_0_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10966_ _06314_ _06921_ _07107_ vssd1 vssd1 vccd1 vccd1 _07306_ sky130_fd_sc_hd__a21bo_1
XANTENNA__09484__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10729__B _06928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12705_ net2265 net258 net385 vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__mux2_1
X_16473_ clknet_leaf_151_wb_clk_i _02227_ _00456_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09302__C net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11291__A2 _06887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13685_ team_01_WB.instance_to_wrap.cpu.c0.count\[12\] _04107_ vssd1 vssd1 vccd1
+ vccd1 _04108_ sky130_fd_sc_hd__and2_1
X_10897_ net520 _06969_ _06970_ _07236_ vssd1 vssd1 vccd1 vccd1 _07237_ sky130_fd_sc_hd__a31o_1
XFILLER_0_26_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10448__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15424_ net1272 vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12636_ net3007 net265 net394 vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09236__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12944__B net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15355_ net1248 vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12567_ net2776 net270 net399 vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__mux2_1
XANTENNA__12436__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14306_ net1324 vssd1 vssd1 vccd1 vccd1 _00100_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11518_ net1550 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[0\] net877 vssd1 vssd1
+ vccd1 vccd1 _03331_ sky130_fd_sc_hd__mux2_1
X_15286_ net1258 vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__inv_2
X_12498_ net3150 net204 net407 vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold208 _02153_ vssd1 vssd1 vccd1 vccd1 net1743 sky130_fd_sc_hd__dlygate4sd3_1
X_17025_ clknet_leaf_55_wb_clk_i _02712_ _01008_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold219 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1754 sky130_fd_sc_hd__dlygate4sd3_1
X_14237_ net1335 vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__inv_2
X_11449_ team_01_WB.instance_to_wrap.cpu.f0.i\[2\] _07672_ net325 vssd1 vssd1 vccd1
+ vccd1 _07749_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13740__A1 net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14168_ _04189_ _04193_ net1823 vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__a21oi_1
X_13119_ net91 net843 net632 net1585 vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__a22o_1
XANTENNA__10480__A _06811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12171__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14099_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[85\] _04245_ _04250_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[125\]
+ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__a22o_1
X_17927_ net1534 vssd1 vssd1 vccd1 vccd1 gpio_oeb[36] sky130_fd_sc_hd__buf_2
Xfanout1270 net1273 vssd1 vssd1 vccd1 vccd1 net1270 sky130_fd_sc_hd__buf_4
X_08660_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[10\] net675 _04981_
+ _04983_ _04987_ vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__a2111o_1
Xfanout1281 net1302 vssd1 vssd1 vccd1 vccd1 net1281 sky130_fd_sc_hd__clkbuf_2
Xfanout1292 net1302 vssd1 vssd1 vccd1 vccd1 net1292 sky130_fd_sc_hd__clkbuf_4
X_17858_ clknet_leaf_125_wb_clk_i team_01_WB.instance_to_wrap.cpu.f0.next_lcd_en _01798_
+ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.SR1.enable sky130_fd_sc_hd__dfrtp_1
XANTENNA__14048__A2 _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16809_ clknet_leaf_40_wb_clk_i _02496_ _00792_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_08591_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[15\] net682 _04928_
+ _04929_ _04930_ vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__a2111o_1
X_17789_ clknet_leaf_95_wb_clk_i net2662 _01729_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11515__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10639__B _06928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09212__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09212_ net1004 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[17\] net887 vssd1
+ vssd1 vccd1 vccd1 _05552_ sky130_fd_sc_hd__and3_1
XANTENNA__13559__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_730 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09143_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[14\] net666 _05457_
+ _05469_ _05477_ vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12346__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09074_ _05405_ _05406_ _05412_ _05413_ vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__or4_1
XANTENNA__12782__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16115__Q team_01_WB.instance_to_wrap.cpu.f0.data_adr\[22\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08025_ team_01_WB.instance_to_wrap.cpu.K0.code\[1\] team_01_WB.instance_to_wrap.cpu.K0.code\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1130_A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold720 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2255 sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2266 sky130_fd_sc_hd__dlygate4sd3_1
Xhold742 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2277 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1228_A net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold753 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2288 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09935__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold764 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2299 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09882__C net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold775 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2310 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout688_A _04773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold786 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[33\] vssd1 vssd1 vccd1 vccd1
+ net2321 sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2332 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12081__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09976_ _06313_ _06315_ vssd1 vssd1 vccd1 vccd1 _06316_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_90_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1016_X net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08927_ net1027 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[6\] net884 vssd1
+ vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__and3_1
XANTENNA__12869__X _03654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout855_A net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout476_X net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1420 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2955 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1431 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2966 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1442 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2977 sky130_fd_sc_hd__dlygate4sd3_1
X_08858_ net1106 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[3\] net931 vssd1
+ vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__and3_1
XANTENNA__14039__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1453 team_01_WB.instance_to_wrap.cpu.f0.num\[7\] vssd1 vssd1 vccd1 vccd1 net2988
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1464 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2999 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1475 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[19\] vssd1 vssd1 vccd1 vccd1
+ net3010 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1486 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net3021 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1497 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3032 sky130_fd_sc_hd__dlygate4sd3_1
X_08789_ net1012 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[0\] net922 vssd1
+ vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout643_X net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10820_ _06967_ _07159_ vssd1 vssd1 vccd1 vccd1 _07160_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_49_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout810_X net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10751_ _06101_ _07089_ _06036_ _06068_ vssd1 vssd1 vccd1 vccd1 _07091_ sky130_fd_sc_hd__a211oi_2
XANTENNA__12470__A1 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_98_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09122__C net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout908_X net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_27_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13470_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] _05592_ vssd1 vssd1
+ vccd1 vccd1 _03931_ sky130_fd_sc_hd__or2_1
XANTENNA__09218__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10682_ _04706_ _05867_ net548 vssd1 vssd1 vccd1 vccd1 _07022_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12421_ net2763 net313 net421 vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12256__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10233__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15140_ net1217 vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12352_ net2183 net309 net428 vssd1 vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11303_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] _05116_ vssd1 vssd1 vccd1
+ vccd1 _07643_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15071_ net1314 vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__inv_2
X_12283_ net1896 net277 net436 vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14022_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[90\] _04240_ _04241_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[90\]
+ vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_112_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11234_ _04738_ _05932_ _06917_ _05707_ _04736_ vssd1 vssd1 vccd1 vccd1 _07574_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__08322__X _04662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_1_0_wb_clk_i_X clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11165_ _06905_ _07254_ _07504_ vssd1 vssd1 vccd1 vccd1 _07505_ sky130_fd_sc_hd__a21oi_1
X_10116_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[6\] net736 _06454_ _06455_
+ vssd1 vssd1 vccd1 vccd1 _06456_ sky130_fd_sc_hd__a211o_1
X_15973_ net1416 vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__inv_2
X_11096_ _07364_ _07379_ _07435_ vssd1 vssd1 vccd1 vccd1 _07436_ sky130_fd_sc_hd__and3b_1
XANTENNA__16686__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11683__X _07884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14924_ net1259 vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__inv_2
X_10047_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[0\] net760 _06380_ _06382_
+ net769 vssd1 vssd1 vccd1 vccd1 _06387_ sky130_fd_sc_hd__a2111o_1
X_17712_ clknet_leaf_125_wb_clk_i _03396_ _01653_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_42_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold80 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 net1615
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 net85 vssd1 vssd1 vccd1 vccd1 net1626 sky130_fd_sc_hd__dlygate4sd3_1
X_14855_ net1390 vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__inv_2
X_17643_ clknet_leaf_157_wb_clk_i _03328_ _01584_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_26_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13806_ team_01_WB.EN_VAL_REG net636 vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__or2_1
X_17574_ clknet_leaf_87_wb_clk_i _03261_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_14786_ net1316 vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__inv_2
X_11998_ net2140 net247 net468 vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__mux2_1
XANTENNA__09457__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16525_ clknet_leaf_157_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[23\]
+ _00508_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13737_ _04511_ _07649_ vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__or2_1
XANTENNA__11264__A2 _07300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10949_ net328 _07288_ _07287_ _07279_ vssd1 vssd1 vccd1 vccd1 _07289_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_27_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_888 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15331__A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16456_ clknet_leaf_8_wb_clk_i _02210_ _00439_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13668_ team_01_WB.instance_to_wrap.a1.curr_state\[0\] _03732_ _04098_ vssd1 vssd1
+ vccd1 vccd1 _04099_ sky130_fd_sc_hd__o21a_1
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15407_ net1296 vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12619_ net3056 net314 net397 vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__mux2_1
XANTENNA__10475__A net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16387_ clknet_leaf_119_wb_clk_i net2859 _00370_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[110\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12166__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13599_ _03907_ _04041_ vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__xnor2_1
X_15338_ net1284 vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15269_ net1286 vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17008_ clknet_leaf_109_wb_clk_i _02695_ _00991_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09917__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09830_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[13\] net790 _06168_
+ _06169_ vssd1 vssd1 vccd1 vccd1 _06170_ sky130_fd_sc_hd__a211o_1
Xfanout507 _06098_ vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__clkbuf_4
Xfanout518 _05260_ vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__clkbuf_2
Xfanout529 net532 vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__clkbuf_4
X_09761_ _06069_ _06100_ vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__and2b_1
XFILLER_0_77_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09207__C net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08712_ net1018 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[5\] net902 vssd1
+ vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__and3_1
X_09692_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] net625 _06030_ _06031_
+ vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__a22o_2
XANTENNA__13492__A3 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08643_ net1020 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[10\] net924 vssd1
+ vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout269_A _07866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08574_ net1000 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[19\] net910
+ vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__and3_1
XANTENNA__09448__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1080_A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10937__X _07277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout436_A net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1178_A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10463__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08781__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12204__A1 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12076__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout603_A _04754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09126_ net1022 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[14\] net903
+ vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_40_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09620__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09057_ net1029 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[12\] net928 vssd1
+ vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_92_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12804__S net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1133_X net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08008_ team_01_WB.instance_to_wrap.cpu.f0.state\[5\] vssd1 vssd1 vccd1 vccd1 _04505_
+ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_145_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_145_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold550 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2085 sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2096 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout972_A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1620_A team_01_WB.instance_to_wrap.cpu.f0.data_adr\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold572 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2107 sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold594 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2129 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout760_X net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09959_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[3\] net789 net775 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06299_ sky130_fd_sc_hd__a22o_1
XANTENNA__09117__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout858_X net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12970_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[116\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[124\]
+ net860 vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__mux2_1
Xhold1250 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2785 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09687__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1261 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2796 sky130_fd_sc_hd__dlygate4sd3_1
X_11921_ net1852 net308 net482 vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__mux2_1
Xhold1272 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2807 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1283 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2818 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12691__A1 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1294 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2829 sky130_fd_sc_hd__dlygate4sd3_1
X_14640_ net1392 vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ net2923 net298 net490 vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__mux2_1
XANTENNA__09439__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10803_ _05657_ net509 vssd1 vssd1 vccd1 vccd1 _07143_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14571_ net1427 vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__inv_2
XANTENNA__11246__A2 _07528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11783_ net1799 net277 net498 vssd1 vssd1 vccd1 vccd1 _03190_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16310_ clknet_leaf_93_wb_clk_i net2206 _00293_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[33\]
+ sky130_fd_sc_hd__dfrtp_1
X_13522_ net198 net194 _07841_ net644 vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__o211a_1
X_10734_ _06912_ _07073_ vssd1 vssd1 vccd1 vccd1 _07074_ sky130_fd_sc_hd__nor2_1
X_17290_ clknet_leaf_31_wb_clk_i _02977_ _01273_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10566__Y _06906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_858 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16241_ clknet_leaf_141_wb_clk_i net1687 _00229_ vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__dfrtp_1
X_13453_ _03900_ _03909_ _03913_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__o21ai_1
X_10665_ net547 _06280_ vssd1 vssd1 vccd1 vccd1 _07005_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_153_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12404_ net2368 net235 net419 vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_153_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16172_ clknet_leaf_1_wb_clk_i _01932_ _00160_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13384_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] _05757_ vssd1 vssd1
+ vccd1 vccd1 _03845_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10757__A1 _04844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10596_ net373 net341 net546 vssd1 vssd1 vccd1 vccd1 _06936_ sky130_fd_sc_hd__mux2_1
XANTENNA__09611__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15123_ net1392 vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__inv_2
XANTENNA__11678__X _07880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12335_ net2394 net242 net429 vssd1 vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__mux2_1
XANTENNA__12714__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15054_ net1297 vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_110_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12266_ net2904 net275 net437 vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__mux2_1
XANTENNA__11706__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14005_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[33\] _04221_ _04252_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[105\]
+ vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__a22o_1
X_11217_ _06814_ _06821_ _07555_ vssd1 vssd1 vccd1 vccd1 _07557_ sky130_fd_sc_hd__or3_1
X_12197_ net1919 net206 net445 vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__mux2_1
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__buf_2
XANTENNA__11182__B2 _06919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__buf_2
X_11148_ net328 _07485_ _07487_ _07478_ vssd1 vssd1 vccd1 vccd1 _07488_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_50_Left_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11079_ net509 _07095_ _05657_ vssd1 vssd1 vccd1 vccd1 _07419_ sky130_fd_sc_hd__and3b_1
XANTENNA__14230__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15956_ net1366 vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_108_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09678__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08866__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14907_ net1247 vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__inv_2
XANTENNA__11573__B team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15887_ net1411 vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08350__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17626_ clknet_leaf_3_wb_clk_i _03311_ _01567_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_14838_ net1258 vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14769_ net1422 vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__inv_2
X_17557_ clknet_leaf_109_wb_clk_i _03244_ _01540_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16508_ clknet_leaf_2_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[6\]
+ _00491_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_08290_ net992 net984 vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__and2_1
X_17488_ clknet_leaf_148_wb_clk_i _03175_ _01471_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09697__C net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10996__A1 _06398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16439_ clknet_leaf_74_wb_clk_i _02193_ _00422_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10748__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12624__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10652__B net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13162__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout315 net316 vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__clkbuf_2
Xfanout326 _07698_ vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__dlymetal6s2s_1
X_09813_ _06138_ _06150_ _06151_ _06152_ vssd1 vssd1 vccd1 vccd1 _06153_ sky130_fd_sc_hd__or4_1
Xfanout337 _06911_ vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__buf_2
Xfanout348 net349 vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__buf_2
XFILLER_0_94_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout359 _03655_ vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10920__A1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout386_A _03570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10920__B2 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09744_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[20\] net821 net755 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _06084_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08877__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09675_ net994 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[22\] net958 vssd1
+ vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout553_A net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1295_A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08626_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[11\] net698 net671 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[11\]
+ _04965_ vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout720_A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08557_ net1078 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[19\] net887
+ vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout341_X net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13622__B1 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout439_X net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout818_A _04634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1083_X net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08488_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[23\] net679 _04818_
+ _04761_ _04786_ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09841__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1250_X net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout606_X net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10450_ net1147 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[26\] net979 vssd1
+ vssd1 vccd1 vccd1 _06790_ sky130_fd_sc_hd__and3b_1
XFILLER_0_150_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09109_ _05445_ _05446_ _05447_ _05448_ vssd1 vssd1 vccd1 vccd1 _05449_ sky130_fd_sc_hd__or4_1
XFILLER_0_21_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10381_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[16\] net786 _06719_
+ _06720_ vssd1 vssd1 vccd1 vccd1 _06721_ sky130_fd_sc_hd__a211o_1
XANTENNA__12534__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12120_ net3100 net307 net458 vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_107_Left_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout975_X net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12051_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[6\] net299 net466 vssd1
+ vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__mux2_1
XANTENNA__13153__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold380 net109 vssd1 vssd1 vccd1 vccd1 net1915 sky130_fd_sc_hd__dlygate4sd3_1
Xhold391 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net1926 sky130_fd_sc_hd__dlygate4sd3_1
X_11002_ _05758_ net504 vssd1 vssd1 vccd1 vccd1 _07342_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_59_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_102_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout860 net867 vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__buf_2
X_15810_ net1200 vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__inv_2
Xfanout871 net872 vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08580__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout882 net883 vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__buf_4
X_16790_ clknet_leaf_29_wb_clk_i _02477_ _00773_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout893 net895 vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__buf_4
XANTENNA__08686__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15741_ net1313 vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__inv_2
X_12953_ net3133 net870 net357 _03711_ vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__a22o_1
XANTENNA__12664__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08868__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1080 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2615 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1091 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2626 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_66_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11904_ net2041 net271 net479 vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_42_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_116_Left_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15672_ net1212 vssd1 vssd1 vccd1 vccd1 _01466_ sky130_fd_sc_hd__inv_2
X_12884_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[27\] _03663_ net1040 vssd1
+ vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__mux2_1
XANTENNA__08983__A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ net1335 vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__inv_2
X_17411_ clknet_leaf_23_wb_clk_i _03098_ _01394_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11835_ net2402 _07855_ net488 vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__mux2_1
XANTENNA__12709__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ clknet_leaf_80_wb_clk_i _03029_ _01325_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09150__Y _05490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10427__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ net1365 vssd1 vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__inv_2
X_11766_ net2759 net274 net496 vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__mux2_1
XANTENNA__10978__A1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09832__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13505_ _03949_ _03963_ vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17273_ clknet_leaf_103_wb_clk_i _02960_ _01256_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10717_ _05902_ _06824_ vssd1 vssd1 vccd1 vccd1 _07057_ sky130_fd_sc_hd__nand2_1
X_14485_ net1411 vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__inv_2
X_11697_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] _07805_ vssd1 vssd1
+ vccd1 vccd1 _07895_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16224_ clknet_leaf_141_wb_clk_i _01984_ _00212_ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13436_ _03890_ _03893_ vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__nor2_1
X_10648_ _06984_ _06987_ net515 vssd1 vssd1 vccd1 vccd1 _06988_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16155_ clknet_leaf_134_wb_clk_i _01918_ _00143_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_125_Left_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13367_ net565 team_01_WB.instance_to_wrap.cpu.f0.next_write_i _04486_ vssd1 vssd1
+ vccd1 vccd1 _03836_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_98_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12444__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14225__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10579_ _06910_ _06917_ vssd1 vssd1 vccd1 vccd1 _06919_ sky130_fd_sc_hd__or2_4
XANTENNA__11201__X _07541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15106_ net1320 vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__inv_2
X_12318_ net2612 net295 net434 vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__mux2_1
X_16086_ clknet_leaf_132_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[8\]
+ _00074_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[8\] sky130_fd_sc_hd__dfrtp_1
X_13298_ team_01_WB.instance_to_wrap.cpu.f0.i\[22\] net610 _07710_ vssd1 vssd1 vccd1
+ vccd1 _03782_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15037_ net1311 vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__inv_2
X_12249_ net1902 net300 net440 vssd1 vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09899__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11584__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16988_ clknet_leaf_60_wb_clk_i _02675_ _00971_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_147_Right_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_134_Left_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15939_ net1367 vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09460_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[29\] net686 net668 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[29\]
+ _05783_ vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__a221o_1
X_08411_ net1170 _04718_ vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__nor2_2
X_17609_ clknet_leaf_86_wb_clk_i _03296_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_09391_ net559 _05570_ vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__nor2_1
XANTENNA__12619__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08342_ net992 net963 vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08273_ net3082 net2346 net1046 vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12354__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1043_A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09339__A1 net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16123__Q team_01_WB.instance_to_wrap.cpu.f0.data_adr\[30\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10950__X _07290_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11146__A1 _06920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07972__A team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_121_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08420__X _04760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09890__C net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout670_A _04800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout768_A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout389_X net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07988_ net1071 vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__inv_2
Xfanout189 net191 vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__clkbuf_2
XANTENNA__14096__B1 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09727_ net377 _05619_ _05731_ _05595_ vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__a211o_1
XANTENNA__12877__X _03659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout556_X net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout935_A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09658_ _04844_ _05733_ vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_2_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10121__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09251__X _05591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08609_ _04751_ _04752_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1 vssd1
+ vccd1 vccd1 _04949_ sky130_fd_sc_hd__o21a_1
XFILLER_0_139_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10397__X _06737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout723_X net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12529__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09589_ _05918_ _05920_ _05925_ _05928_ vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__or4_1
XFILLER_0_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11620_ _07820_ _07833_ vssd1 vssd1 vccd1 vccd1 _07834_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_61_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08078__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09814__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10557__B net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_132_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_154_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11551_ net1728 net1173 vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__and2_1
XANTENNA__09130__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10502_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[31\] net745 _06834_ _06838_
+ _06840_ vssd1 vssd1 vccd1 vccd1 _06842_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_150_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14270_ net1225 vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_150_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14020__B1 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11482_ net366 _07768_ net3101 net874 vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_135_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13221_ net2743 net353 net349 team_01_WB.instance_to_wrap.cpu.f0.i\[29\] vssd1 vssd1
+ vccd1 vccd1 _01929_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10433_ _06769_ _06770_ _06771_ _06772_ vssd1 vssd1 vccd1 vccd1 _06773_ sky130_fd_sc_hd__or4_1
XANTENNA__12264__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input64_A wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13152_ net1636 net850 net842 net1589 vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__a22o_1
X_10364_ _06691_ _06692_ _06702_ _06703_ vssd1 vssd1 vccd1 vccd1 _06704_ sky130_fd_sc_hd__or4_1
X_12103_ net2459 net269 net455 vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__mux2_1
XANTENNA__13126__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17960_ net1475 vssd1 vssd1 vccd1 vccd1 la_data_out[2] sky130_fd_sc_hd__buf_2
X_13083_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[3\] net3084 net861 vssd1 vssd1
+ vccd1 vccd1 _02042_ sky130_fd_sc_hd__mux2_1
X_10295_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[19\] net763 net622 vssd1
+ vssd1 vccd1 vccd1 _06635_ sky130_fd_sc_hd__o21a_1
X_16911_ clknet_leaf_31_wb_clk_i _02598_ _00894_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_12034_ net2217 net203 net463 vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_148_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17891_ net1513 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
XFILLER_0_18_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11608__S net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08553__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16842_ clknet_leaf_11_wb_clk_i _02529_ _00825_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10360__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout690 _04772_ vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__clkbuf_8
X_16773_ clknet_leaf_46_wb_clk_i _02460_ _00756_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13985_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[8\] _04226_ _04256_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[40\]
+ _04276_ vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__a221o_1
XFILLER_0_125_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15724_ net1260 vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__inv_2
X_12936_ net357 _03699_ _03700_ net870 net1764 vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__a32o_1
XANTENNA__10112__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12947__B net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15655_ net1390 vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__inv_2
XANTENNA__12439__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12867_ net585 _07756_ vssd1 vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__or2_2
X_11818_ net1905 net292 net494 vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__mux2_1
X_14606_ net1357 vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09266__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15586_ net1319 vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__inv_2
X_12798_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[10\] _07531_ net1035 vssd1 vssd1
+ vccd1 vccd1 _03627_ sky130_fd_sc_hd__mux2_1
XANTENNA__09805__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16208__Q net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14537_ net1364 vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17325_ clknet_leaf_68_wb_clk_i _03012_ _01308_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11749_ _04501_ _07936_ net615 vssd1 vssd1 vccd1 vccd1 _07937_ sky130_fd_sc_hd__mux2_4
XFILLER_0_44_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17256_ clknet_leaf_62_wb_clk_i _02943_ _01239_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_14468_ net1356 vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__inv_2
XANTENNA__14011__B1 _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13419_ _03877_ _03878_ _03869_ vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__a21o_1
X_16207_ clknet_leaf_124_wb_clk_i _01967_ _00195_ vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17187_ clknet_leaf_25_wb_clk_i _02874_ _01170_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12174__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14399_ net1307 vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__inv_2
XANTENNA__10179__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16138_ clknet_leaf_128_wb_clk_i _01901_ _00126_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08792__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08960_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[6\] net704 _05296_ _05299_
+ vssd1 vssd1 vccd1 vccd1 _05300_ sky130_fd_sc_hd__o22a_4
XFILLER_0_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16069_ clknet_leaf_156_wb_clk_i _01862_ _00057_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\]
+ sky130_fd_sc_hd__dfstp_4
XANTENNA__10770__X _07110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11128__B2 _06906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13522__C1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08891_ net1025 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[2\] net919 vssd1
+ vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__and3_1
XANTENNA__11518__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_75 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14078__B1 _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10351__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09512_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[29\] net761 net751 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[29\]
+ _05850_ vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__a221o_1
XANTENNA__11300__A1 _05153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09443_ net1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[29\] net903
+ vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__and3_1
XANTENNA__12349__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout251_A _07904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09257__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09374_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[26\] net692 net659 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08325_ net1165 net1166 net1158 net1162 vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__and4b_1
XFILLER_0_145_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12800__B2 _03628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1258_A net1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08256_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[25\] net2429 net1056 vssd1 vssd1
+ vccd1 vccd1 _03431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14002__B1 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09885__C net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12084__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08187_ net2730 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[86\] net1044 vssd1 vssd1
+ vccd1 vccd1 _03500_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1425_A net1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout885_A net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08798__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11119__A1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10080_ net1138 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[7\] net975 vssd1
+ vssd1 vccd1 vccd1 _06420_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout673_X net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_6_0_wb_clk_i_X clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08535__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14069__B1 _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09125__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout938_X net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13770_ team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[3\] _04146_ vssd1 vssd1
+ vccd1 vccd1 _04157_ sky130_fd_sc_hd__or2_1
X_10982_ net558 _07311_ _07321_ net328 vssd1 vssd1 vccd1 vccd1 _07322_ sky130_fd_sc_hd__a22o_1
XANTENNA__08964__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12721_ team_01_WB.instance_to_wrap.a1.WRITE_I team_01_WB.instance_to_wrap.cpu.RU0.state\[1\]
+ _03571_ vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__or3_4
XFILLER_0_69_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12259__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11163__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15440_ net1276 vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12652_ net2893 net314 net392 vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09248__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11603_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\]
+ _07819_ vssd1 vssd1 vccd1 vccd1 _07820_ sky130_fd_sc_hd__and3_2
XFILLER_0_33_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15371_ net1396 vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12583_ net1866 net309 net400 vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__mux2_1
X_14322_ net1330 vssd1 vssd1 vccd1 vccd1 _00116_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17110_ clknet_leaf_12_wb_clk_i _02797_ _01093_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11534_ net2108 net1174 net589 net1134 vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__a22o_1
Xwire321 net322 vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_111_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17041_ clknet_leaf_114_wb_clk_i _02728_ _01024_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11399__A team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14253_ net1226 vssd1 vssd1 vccd1 vccd1 _00047_ sky130_fd_sc_hd__inv_2
X_11465_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[30\] net579 vssd1 vssd1 vccd1
+ vccd1 _07760_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_78_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13204_ net4 net836 net629 net2150 vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__o22a_1
XFILLER_0_150_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10416_ net1132 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[27\] net968
+ vssd1 vssd1 vccd1 vccd1 _06756_ sky130_fd_sc_hd__and3_1
X_14184_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[12\] _04453_ net1427 vssd1
+ vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11396_ _07668_ _07697_ _07699_ _07714_ vssd1 vssd1 vccd1 vccd1 _07721_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_115_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13135_ net1733 net846 net633 team_01_WB.instance_to_wrap.a1.ADR_I\[8\] vssd1 vssd1
+ vccd1 vccd1 _02006_ sky130_fd_sc_hd__a22o_1
XANTENNA__08774__A2 _05110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10347_ net1135 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[17\] net965
+ vssd1 vssd1 vccd1 vccd1 _06687_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17943_ net1458 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
X_13066_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[20\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[28\]
+ net854 vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__mux2_1
X_10278_ net1128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[19\] net970
+ vssd1 vssd1 vccd1 vccd1 _06618_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1430 net38 vssd1 vssd1 vccd1 vccd1 net1430 sky130_fd_sc_hd__buf_4
X_12017_ net1772 net276 net470 vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17874_ clknet_leaf_138_wb_clk_i _03549_ _01814_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11530__B2 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16825_ clknet_leaf_71_wb_clk_i _02512_ _00808_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16756_ clknet_leaf_21_wb_clk_i _02443_ _00739_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13968_ _04225_ _04232_ vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__nor2_4
XANTENNA__10097__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[7\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15707_ net1251 vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__inv_2
X_12919_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[17\] net1040 vssd1 vssd1 vccd1
+ vccd1 _03689_ sky130_fd_sc_hd__or2_1
XANTENNA__12169__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13899_ net571 _04200_ _04201_ vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__and3_1
X_16687_ clknet_leaf_33_wb_clk_i _02374_ _00670_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15638_ net1247 vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09239__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15569_ net1420 vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11801__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08110_ net1070 team_01_WB.instance_to_wrap.cpu.f0.num\[8\] vssd1 vssd1 vccd1 vccd1
+ _04580_ sky130_fd_sc_hd__nor2_1
X_17308_ clknet_leaf_59_wb_clk_i _02995_ _01291_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09090_ net1011 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[13\] net887 vssd1
+ vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__and3_1
X_08041_ net1670 net568 net346 team_01_WB.instance_to_wrap.cpu.f0.i\[14\] vssd1 vssd1
+ vccd1 vccd1 _03550_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17239_ clknet_leaf_13_wb_clk_i _02926_ _01222_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold902 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold913 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[82\] vssd1 vssd1 vccd1 vccd1
+ net2448 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap621 _04730_ vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_842 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold924 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2459 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold935 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold946 _02090_ vssd1 vssd1 vccd1 vccd1 net2481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2492 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08765__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold968 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2503 sky130_fd_sc_hd__dlygate4sd3_1
X_09992_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[2\] net735 _06330_ _06331_
+ vssd1 vssd1 vccd1 vccd1 _06332_ sky130_fd_sc_hd__a211o_1
XANTENNA__12632__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold979 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2514 sky130_fd_sc_hd__dlygate4sd3_1
X_08943_ net1111 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[6\] net907 vssd1
+ vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_32_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout299_A _07921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1602 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net3137 sky130_fd_sc_hd__dlygate4sd3_1
X_08874_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[3\] net694 net682 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[3\]
+ _05204_ vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_4_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1613 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net3148 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1006_A net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1624 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net3159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1635 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1646 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 net3181
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout466_A _07954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09478__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08308__B_N net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12079__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout633_A _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09426_ net1097 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[28\] net909
+ net650 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[28\] vssd1 vssd1 vccd1
+ vccd1 _05766_ sky130_fd_sc_hd__a32o_1
XFILLER_0_137_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12874__Y _03657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09357_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[25\] net691 net663 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout800_A net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10675__X _07015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout421_X net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1163_X net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12785__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08308_ net1162 net1168 net1164 net1158 vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__and4bb_2
X_09288_ net1009 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[22\] net878
+ vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__and3_1
XFILLER_0_62_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08239_ net2372 net2440 net1053 vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1428_X net1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11250_ _05967_ _06748_ _06749_ vssd1 vssd1 vccd1 vccd1 _07590_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_95_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09402__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout790_X net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout888_X net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10201_ net1140 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[8\] net975 vssd1
+ vssd1 vccd1 vccd1 _06541_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12542__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11181_ _06532_ _07190_ net343 vssd1 vssd1 vccd1 vccd1 _07521_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10132_ _06442_ _06471_ _06470_ vssd1 vssd1 vccd1 vccd1 _06472_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_73_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10570__B _04738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10063_ _06339_ _06342_ vssd1 vssd1 vccd1 vccd1 _06403_ sky130_fd_sc_hd__xnor2_1
X_14940_ net1244 vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__inv_2
XANTENNA__11512__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input27_A DAT_I[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14871_ net1213 vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_141_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16610_ clknet_leaf_77_wb_clk_i _02297_ _00593_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11682__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13822_ net1701 net832 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[15\]
+ sky130_fd_sc_hd__and2_1
X_17590_ clknet_leaf_130_wb_clk_i _03277_ _01549_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.code\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13265__B2 _04621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13753_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[9\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[11\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[10\] vssd1 vssd1 vccd1 vccd1 _04142_
+ sky130_fd_sc_hd__and3_1
X_16541_ clknet_leaf_6_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[7\]
+ _00524_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_10965_ _05263_ _07303_ _07304_ vssd1 vssd1 vccd1 vccd1 _07305_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_70_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12704_ net1867 net231 net385 vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13684_ team_01_WB.instance_to_wrap.cpu.c0.count\[10\] team_01_WB.instance_to_wrap.cpu.c0.count\[11\]
+ _04106_ vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__and3_1
X_16472_ clknet_leaf_141_wb_clk_i _02226_ _00455_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10896_ net520 _07138_ vssd1 vssd1 vccd1 vccd1 _07236_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15423_ net1319 vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__inv_2
X_12635_ net1946 net233 net391 vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12717__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11621__S net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13402__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15354_ net1372 vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12566_ net2863 net241 net401 vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__mux2_1
XANTENNA__09641__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08995__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14305_ net1324 vssd1 vssd1 vccd1 vccd1 _00099_ sky130_fd_sc_hd__inv_2
X_11517_ net1551 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[1\] net877 vssd1 vssd1
+ vccd1 vccd1 _03332_ sky130_fd_sc_hd__mux2_1
X_15285_ net1287 vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12497_ net2997 net273 net409 vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17024_ clknet_leaf_45_wb_clk_i _02711_ _01007_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold209 team_01_WB.instance_to_wrap.cpu.f0.write_data\[19\] vssd1 vssd1 vccd1 vccd1
+ net1744 sky130_fd_sc_hd__dlygate4sd3_1
X_14236_ net1335 vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11448_ _07674_ _07748_ vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__nor2_1
X_14167_ _04189_ _04193_ _04444_ net1426 vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__a211oi_1
XANTENNA__12452__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13740__A2 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11379_ _07707_ vssd1 vssd1 vccd1 vccd1 _07708_ sky130_fd_sc_hd__inv_2
XANTENNA__10761__A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11751__A1 _07476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13118_ net92 net844 net633 net1559 vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__a22o_1
X_14098_ _04378_ _04380_ _04382_ _04384_ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__or4_1
X_17926_ net1533 vssd1 vssd1 vccd1 vccd1 gpio_oeb[35] sky130_fd_sc_hd__buf_2
X_13049_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[37\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[45\]
+ net859 vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1260 net1269 vssd1 vssd1 vccd1 vccd1 net1260 sky130_fd_sc_hd__buf_4
XANTENNA__17240__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1271 net1273 vssd1 vssd1 vccd1 vccd1 net1271 sky130_fd_sc_hd__buf_2
Xfanout1282 net1285 vssd1 vssd1 vccd1 vccd1 net1282 sky130_fd_sc_hd__buf_4
X_17857_ clknet_leaf_121_wb_clk_i net1760 _01797_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[127\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1293 net1301 vssd1 vssd1 vccd1 vccd1 net1293 sky130_fd_sc_hd__buf_4
XANTENNA__11592__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15064__A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16808_ clknet_leaf_63_wb_clk_i _02495_ _00791_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_08590_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[15\] net673 net657 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__a22o_1
X_17788_ clknet_leaf_91_wb_clk_i net2762 _01728_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16739_ clknet_leaf_26_wb_clk_i _02426_ _00722_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09211_ net1087 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[17\] net896
+ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12627__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12767__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09142_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[14\] _04789_ _05463_
+ _05465_ _05476_ vssd1 vssd1 vccd1 vccd1 _05482_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_8_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09073_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[12\] net675 _05383_
+ _05386_ _05394_ vssd1 vssd1 vccd1 vccd1 _05413_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_20_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16045__D net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout214_A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08024_ team_01_WB.instance_to_wrap.cpu.f0.state\[5\] _04506_ _04511_ net586 _04519_
+ vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_130_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold710 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2245 sky130_fd_sc_hd__dlygate4sd3_1
Xhold721 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2256 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold732 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2267 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13192__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold743 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2278 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold754 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2289 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12362__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold765 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2300 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1123_A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold776 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2311 sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 _03439_ vssd1 vssd1 vccd1 vccd1 net2322 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08779__C net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09975_ net527 _06282_ _06314_ net377 vssd1 vssd1 vccd1 vccd1 _06315_ sky130_fd_sc_hd__a22o_1
Xhold798 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2333 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08926_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] net597 net596 vssd1 vssd1
+ vccd1 vccd1 _05266_ sky130_fd_sc_hd__and3_1
Xhold1410 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[64\] vssd1 vssd1 vccd1 vccd1
+ net2945 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07980__A team_01_WB.instance_to_wrap.cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09163__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1421 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[96\] vssd1 vssd1 vccd1 vccd1
+ net2956 sky130_fd_sc_hd__dlygate4sd3_1
X_08857_ net1102 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[3\] net915 vssd1
+ vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__and3_1
Xhold1432 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2967 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout750_A _04680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout371_X net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1443 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2978 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1454 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2989 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout469_X net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1465 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[81\] vssd1 vssd1 vccd1 vccd1
+ net3000 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout848_A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08910__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1476 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net3011 sky130_fd_sc_hd__dlygate4sd3_1
X_08788_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[0\] net695 _05125_ _05126_
+ _05127_ vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__a2111o_1
Xhold1487 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3022 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13247__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold1498 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[22\] vssd1 vssd1 vccd1 vccd1
+ net3033 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10750_ _06101_ _07089_ _06068_ vssd1 vssd1 vccd1 vccd1 _07090_ sky130_fd_sc_hd__a21o_1
XANTENNA__09871__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_958 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09409_ _05742_ _05744_ _05746_ _05748_ vssd1 vssd1 vccd1 vccd1 _05749_ sky130_fd_sc_hd__or4_1
XANTENNA__09700__A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout803_X net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12537__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10681_ _05901_ _06825_ _06827_ net343 vssd1 vssd1 vccd1 vccd1 _07021_ sky130_fd_sc_hd__a31o_1
XANTENNA__12758__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12420_ net2356 net320 net422 vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09623__B1 _05961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10565__B net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12351_ net2666 net292 net429 vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_67_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_134_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11302_ _07640_ _07641_ vssd1 vssd1 vccd1 vccd1 _07642_ sky130_fd_sc_hd__and2b_1
XFILLER_0_22_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15070_ net1350 vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__inv_2
X_12282_ net2410 net301 net436 vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14021_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[42\] _04256_ _04264_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[106\]
+ vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11677__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11233_ _06966_ _07265_ vssd1 vssd1 vccd1 vccd1 _07573_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_112_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10581__A _04710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12272__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10536__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08689__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12930__B1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11164_ _05262_ _07467_ _07503_ net531 vssd1 vssd1 vccd1 vccd1 _07504_ sky130_fd_sc_hd__a22o_1
X_10115_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[6\] _04636_ net784 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06455_ sky130_fd_sc_hd__a22o_1
X_11095_ _07334_ _07391_ _07398_ _07434_ vssd1 vssd1 vccd1 vccd1 _07435_ sky130_fd_sc_hd__and4b_1
X_15972_ net1366 vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__inv_2
X_17711_ clknet_leaf_125_wb_clk_i _03395_ _01652_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14923_ net1424 vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__inv_2
X_10046_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[0\] net756 _06370_ _06377_
+ _06381_ vssd1 vssd1 vccd1 vccd1 _06386_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_136_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold70 _02019_ vssd1 vssd1 vccd1 vccd1 net1605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 net128 vssd1 vssd1 vccd1 vccd1 net1616 sky130_fd_sc_hd__dlygate4sd3_1
X_17642_ clknet_leaf_157_wb_clk_i _03327_ _01583_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold92 _02017_ vssd1 vssd1 vccd1 vccd1 net1627 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_69_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14854_ net1400 vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__inv_2
X_13805_ _04159_ _04181_ _04183_ vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__a21bo_1
X_17573_ clknet_leaf_87_wb_clk_i _03260_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_14785_ net1240 vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__inv_2
X_11997_ net2964 net211 net467 vssd1 vssd1 vccd1 vccd1 _02986_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16524_ clknet_leaf_159_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[22\]
+ _00507_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15612__A net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10948_ _07283_ _07286_ net526 vssd1 vssd1 vccd1 vccd1 _07288_ sky130_fd_sc_hd__mux2_1
X_13736_ team_01_WB.instance_to_wrap.cpu.K0.keyvalid net1700 _04523_ _04135_ vssd1
+ vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__a31o_1
XANTENNA__09862__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16455_ clknet_leaf_31_wb_clk_i _02209_ _00438_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12447__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10756__A net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13667_ net3153 _04097_ vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__nand2_1
X_10879_ _07028_ _07036_ net519 vssd1 vssd1 vccd1 vccd1 _07219_ sky130_fd_sc_hd__mux2_1
XANTENNA__14228__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12749__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15406_ net1297 vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12618_ net2933 net318 net398 vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__mux2_1
X_16386_ clknet_leaf_92_wb_clk_i _02140_ _00369_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[109\]
+ sky130_fd_sc_hd__dfstp_1
X_13598_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] _05381_ _04029_ vssd1
+ vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09614__B1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15337_ net1293 vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__inv_2
X_12549_ net2671 net293 net405 vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11972__A1 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_1 _03570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15268_ net1219 vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__inv_2
X_17007_ clknet_leaf_31_wb_clk_i _02694_ _00990_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12182__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14219_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[13\] vssd1 vssd1 vccd1
+ vccd1 _02268_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10491__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15199_ net1313 vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__inv_2
XANTENNA__10527__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11724__B2 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout508 _06065_ vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout519 net520 vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__clkbuf_4
X_09760_ _06099_ net507 vssd1 vssd1 vccd1 vccd1 _06100_ sky130_fd_sc_hd__nand2b_1
X_08711_ net1018 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[5\] net885 vssd1
+ vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__and3_1
XANTENNA__09145__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17909_ net1520 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
X_09691_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[22\] net763 net622 vssd1
+ vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__o21a_1
Xfanout1090 net1096 vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__buf_2
X_08642_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[10\] net941
+ vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__and3_1
XFILLER_0_83_75 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08573_ net1000 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[19\] net918 vssd1
+ vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1073_A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout429_A _07965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09125_ net1110 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[14\] net927
+ vssd1 vssd1 vccd1 vccd1 _05465_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout217_X net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1338_A net1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09056_ net1029 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[12\] net894
+ vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_92_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09893__C net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout798_A net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08007_ net1175 vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__clkinv_4
XANTENNA__13165__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold540 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2075 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12092__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold551 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[3\] vssd1 vssd1 vccd1 vccd1
+ net2086 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11715__A1 _07290_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12912__B1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold562 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2097 sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[19\] vssd1 vssd1 vccd1 vccd1
+ net2108 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09384__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_49_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_12_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold584 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[30\] vssd1 vssd1 vccd1 vccd1 net2119
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2130 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08302__C net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08592__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09958_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[3\] net737 _06291_ _06295_
+ _06297_ vssd1 vssd1 vccd1 vccd1 _06298_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_95_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08909_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[2\] net668 _05231_ _05235_
+ _05237_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout753_X net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09889_ net1157 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[5\] net946 vssd1
+ vssd1 vccd1 vccd1 _06229_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_114_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_114_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold1240 _03453_ vssd1 vssd1 vccd1 vccd1 net2775 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13217__A net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1251 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2786 sky130_fd_sc_hd__dlygate4sd3_1
X_11920_ net2069 net311 net480 vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__mux2_1
Xhold1262 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[30\] vssd1 vssd1 vccd1 vccd1
+ net2797 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1273 team_01_WB.instance_to_wrap.cpu.f0.num\[24\] vssd1 vssd1 vccd1 vccd1 net2808
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10151__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1284 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2819 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1295 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2830 sky130_fd_sc_hd__dlygate4sd3_1
X_11851_ net2562 net279 net488 vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__mux2_1
XANTENNA__09133__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout920_X net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10802_ _05657_ net509 vssd1 vssd1 vccd1 vccd1 _07142_ sky130_fd_sc_hd__or2_1
XANTENNA__10279__C net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14570_ net1366 vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__inv_2
X_11782_ net1868 net303 net495 vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__mux2_1
XANTENNA__09844__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13640__A1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10847__Y _07187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08972__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10733_ _05781_ _05898_ vssd1 vssd1 vccd1 vccd1 _07073_ sky130_fd_sc_hd__and2_1
X_13521_ _03944_ _03976_ vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_24_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12267__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16240_ clknet_leaf_140_wb_clk_i net1645 _00228_ vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__dfrtp_1
X_13452_ _03904_ _03906_ _03912_ _03911_ vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__a31oi_1
X_10664_ _07000_ _07003_ net517 vssd1 vssd1 vccd1 vccd1 _07004_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12403_ net2969 net240 net419 vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11959__X _07952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13383_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] _05780_ vssd1 vssd1
+ vccd1 vccd1 _03844_ sky130_fd_sc_hd__xor2_1
X_16171_ clknet_leaf_3_wb_clk_i _00013_ _00159_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_153_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_88_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10595_ net553 _06902_ vssd1 vssd1 vccd1 vccd1 _06935_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10757__A2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15122_ net1291 vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__inv_2
X_12334_ net2065 _07858_ net428 vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__mux2_1
XANTENNA__13156__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15053_ net1267 vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12265_ net3013 net207 net437 vssd1 vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11706__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10509__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14004_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[9\] _04253_ _04266_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12903__B1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11216_ _06814_ _07555_ _06821_ vssd1 vssd1 vccd1 vccd1 _07556_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09375__A2 _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12196_ net1979 net246 net445 vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__mux2_1
XANTENNA__11182__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__buf_2
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 ADR_O[26] sky130_fd_sc_hd__buf_2
X_11147_ _06906_ _07319_ _07483_ net526 vssd1 vssd1 vccd1 vccd1 _07487_ sky130_fd_sc_hd__o22a_1
XANTENNA__09605__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14120__A2 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11078_ _07415_ _07416_ _07417_ _07357_ vssd1 vssd1 vccd1 vccd1 _07418_ sky130_fd_sc_hd__o31a_1
X_15955_ net1367 vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__inv_2
XANTENNA__10250__S net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10029_ _06366_ _06367_ _06368_ vssd1 vssd1 vccd1 vccd1 _06369_ sky130_fd_sc_hd__and3_1
X_14906_ net1371 vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__inv_2
X_15886_ net1408 vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10142__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17625_ clknet_leaf_5_wb_clk_i net1806 _01566_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_14837_ net1275 vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__inv_2
XANTENNA__09043__C net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12966__A net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17556_ clknet_leaf_67_wb_clk_i _03243_ _01539_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09835__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12877__B1_N net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14768_ net1278 vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__inv_2
XANTENNA__09978__C net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09340__A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16507_ clknet_leaf_2_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[5\]
+ _00490_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13719_ team_01_WB.instance_to_wrap.cpu.c0.count\[10\] _04106_ net3151 vssd1 vssd1
+ vccd1 vccd1 _04129_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12177__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17487_ clknet_leaf_34_wb_clk_i _03174_ _01470_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14699_ net1210 vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__inv_2
XANTENNA__10996__A2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16438_ clknet_leaf_71_wb_clk_i _02192_ _00421_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12905__S net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16369_ clknet_leaf_99_wb_clk_i _02123_ _00352_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[92\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_147_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08810__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13147__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout305 _07935_ vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__buf_2
XANTENNA__10905__C1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11173__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout316 _07939_ vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__dlymetal6s2s_1
X_09812_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[14\] net822 net798 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06152_ sky130_fd_sc_hd__a22o_1
Xfanout327 _07101_ vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__buf_2
XANTENNA__12640__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout338 _06903_ vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__clkbuf_4
Xfanout349 _03742_ vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__buf_2
XFILLER_0_94_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09743_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[20\] net777 net746 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__a22o_1
XANTENNA__14111__A2 _04244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout281_A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_A net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11109__X _07449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09674_ net994 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[22\] net972 vssd1
+ vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__and3_1
X_08625_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[11\] net693 net674 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08629__A1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08556_ net1077 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[19\] net918
+ vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__and3_1
XANTENNA__13622__A1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09888__C net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11633__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_122_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12087__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1396_A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[23\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08487_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[23\] net693 _04774_ _04781_
+ _04826_ vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout713_A net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout334_X net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1076_X net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout501_X net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09108_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[13\] net656 _05420_
+ _05426_ _05439_ vssd1 vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_131_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10380_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[16\] net784 net745 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06720_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13994__X _04286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09039_ _05264_ _05265_ _05302_ _05377_ vssd1 vssd1 vccd1 vccd1 _05379_ sky130_fd_sc_hd__or4b_2
X_12050_ net2870 net277 net464 vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__mux2_1
XANTENNA__09357__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold370 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1905 sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 _01976_ vssd1 vssd1 vccd1 vccd1 net1916 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09128__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11001_ _07072_ _07073_ _07340_ _07045_ vssd1 vssd1 vccd1 vccd1 _07341_ sky130_fd_sc_hd__o211ai_2
XANTENNA_fanout968_X net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08565__B1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold392 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1927 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12550__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15427__A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout850 net851 vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__clkbuf_4
Xfanout861 net867 vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14102__A2 _04241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout872 net873 vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__clkbuf_4
Xfanout883 _04803_ vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__clkbuf_4
Xfanout894 net895 vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__clkbuf_4
X_15740_ net1245 vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__inv_2
X_12952_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[6\] _05300_ net1039 vssd1
+ vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__mux2_1
XANTENNA__10124__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1070 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2605 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1081 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[48\] vssd1 vssd1 vccd1 vccd1
+ net2616 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1092 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[18\] vssd1 vssd1 vccd1 vccd1
+ net2627 sky130_fd_sc_hd__dlygate4sd3_1
X_11903_ net2754 net241 net481 vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__mux2_1
X_15671_ net1214 vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__inv_2
X_12883_ _05756_ net578 net361 vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__o21ba_2
X_17410_ clknet_leaf_76_wb_clk_i _03097_ _01393_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ net1305 vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ net2357 net274 net489 vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__mux2_1
XANTENNA__13613__A1 team_01_WB.instance_to_wrap.cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09160__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17341_ clknet_leaf_75_wb_clk_i _03028_ _01324_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11765_ net3037 net208 net496 vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__mux2_1
X_14553_ net1411 vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_155_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_82_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_56_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10716_ _07020_ _07021_ _07053_ vssd1 vssd1 vccd1 vccd1 _07056_ sky130_fd_sc_hd__o21ai_4
X_13504_ _03842_ _03843_ vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__and2_1
X_17272_ clknet_leaf_49_wb_clk_i _02959_ _01255_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14484_ net1406 vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__inv_2
X_11696_ net718 _07520_ net616 _07893_ vssd1 vssd1 vccd1 vccd1 _07894_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_11_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16223_ clknet_leaf_135_wb_clk_i _01983_ _00211_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10647_ _06985_ _06986_ net536 vssd1 vssd1 vccd1 vccd1 _06987_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13435_ _03889_ _03892_ _03895_ vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__or3_1
XANTENNA__13410__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16154_ clknet_leaf_137_wb_clk_i _01917_ _00142_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13366_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[10\] _03835_ net827 vssd1 vssd1
+ vccd1 vccd1 _01878_ sky130_fd_sc_hd__mux2_1
X_10578_ _06910_ _06917_ vssd1 vssd1 vccd1 vccd1 _06918_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13129__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15105_ net1239 vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__inv_2
X_12317_ net2519 net298 net434 vssd1 vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__mux2_1
X_16085_ clknet_leaf_132_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[7\]
+ _00073_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[7\] sky130_fd_sc_hd__dfrtp_1
X_13297_ net586 _07649_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.next_write_i
+ sky130_fd_sc_hd__or2_1
XANTENNA__08998__X _05338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09348__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12248_ net2937 net282 net442 vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__mux2_1
X_15036_ net1246 vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12179_ net1871 net250 net450 vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__mux2_1
XANTENNA__12460__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10363__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14241__A net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16987_ clknet_leaf_71_wb_clk_i _02674_ _00970_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15938_ net1363 vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__inv_2
XANTENNA__10115__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15869_ net1203 vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__inv_2
XANTENNA__13144__X _03734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08410_ _04736_ net563 vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__nand2_2
XANTENNA__11804__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17608_ clknet_leaf_86_wb_clk_i _03295_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09390_ net376 net342 _05493_ net559 vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__a31o_1
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08341_ net1133 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[30\] net951
+ vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__and3_1
X_17539_ clknet_leaf_26_wb_clk_i _03226_ _01522_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09501__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08272_ net2328 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[1\] net1056 vssd1 vssd1
+ vccd1 vccd1 _03415_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13368__B1 _07650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12635__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09587__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08414__A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_726 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09229__B _04919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10155__S net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1036_A net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout496_A net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12370__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1203_A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08787__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input1_A ACK_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07987_ net1070 vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout663_A _04806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09726_ _05570_ _05618_ _05594_ net559 vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__a211o_1
XANTENNA__10106__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09511__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09657_ net510 vssd1 vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_2_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout830_A net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout451_X net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11714__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08608_ _04947_ vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__inv_2
X_09588_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[25\] net789 net770 _05926_
+ _05927_ vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_132_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08539_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[18\] net676 _04856_
+ _04865_ _04870_ vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_132_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11082__A1 _04844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11550_ net2082 net1173 vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__and2_1
XFILLER_0_135_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13359__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10501_ net1130 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[31\] net970
+ vssd1 vssd1 vccd1 vccd1 _06841_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12545__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11481_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[22\] net579 vssd1 vssd1 vccd1
+ vccd1 _07768_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_150_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10854__A net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13220_ net2669 net355 net351 team_01_WB.instance_to_wrap.cpu.f0.i\[30\] vssd1 vssd1
+ vccd1 vccd1 _01930_ sky130_fd_sc_hd__a22o_1
X_10432_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[27\] net791 net779 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06772_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_862 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08324__A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10573__B _04743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13151_ net125 net849 net841 net2197 vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10363_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[17\] net786 net748 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _06703_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_59_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12102_ net2245 net243 net457 vssd1 vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13082_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[4\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[12\]
+ net854 vssd1 vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__mux2_1
XANTENNA_input57_A wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10294_ _06621_ _06626_ _06633_ vssd1 vssd1 vccd1 vccd1 _06634_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_76_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12334__A1 _07858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16910_ clknet_leaf_27_wb_clk_i _02597_ _00893_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13531__B1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12033_ net2315 net273 net465 vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__mux2_1
XANTENNA__12280__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17890_ net107 vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_148_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12885__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16841_ clknet_leaf_40_wb_clk_i _02528_ _00824_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09750__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout680 _04787_ vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__buf_6
Xfanout691 _04772_ vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__clkbuf_8
X_16772_ clknet_leaf_82_wb_clk_i _02459_ _00755_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08994__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13984_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[32\] _04230_ _04258_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[56\]
+ vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15723_ net1396 vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__inv_2
X_12935_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[12\] net1039 vssd1 vssd1 vccd1
+ vccd1 _03700_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_122_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13405__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15654_ net1384 vssd1 vssd1 vccd1 vccd1 _01448_ sky130_fd_sc_hd__inv_2
X_12866_ net1178 team_01_WB.instance_to_wrap.cpu.RU0.state\[6\] team_01_WB.instance_to_wrap.a1.WRITE_I
+ vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14605_ net1358 vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__inv_2
X_11817_ net2544 net297 net494 vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15585_ net1278 vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__inv_2
X_12797_ net1634 net639 net607 _03626_ vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_859 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17324_ clknet_leaf_20_wb_clk_i _03011_ _01307_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13745__A_N net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14536_ net1352 vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__inv_2
X_11748_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[2\] _07489_ net716 vssd1 vssd1
+ vccd1 vccd1 _07936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17255_ clknet_leaf_100_wb_clk_i _02942_ _01238_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12455__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14467_ net1358 vssd1 vssd1 vccd1 vccd1 _00261_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11679_ net3028 net264 net500 vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__mux2_1
X_16206_ clknet_leaf_124_wb_clk_i net1771 _00194_ vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__dfrtp_1
X_13418_ _03869_ _03878_ vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__nand2b_1
X_17186_ clknet_leaf_55_wb_clk_i _02873_ _01169_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_144_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14398_ net1335 vssd1 vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16137_ clknet_leaf_137_wb_clk_i _01900_ _00125_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13349_ net1671 net827 _03822_ vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16068_ clknet_leaf_156_wb_clk_i _01861_ _00056_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_59_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09726__C1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15019_ net1396 vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__inv_2
X_08890_ net1107 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[2\] net907 vssd1
+ vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__and3_1
XANTENNA__10703__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12876__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08369__A_N team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10004__A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09511_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[29\] net737 _05841_
+ _05842_ _05845_ vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_79_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08701__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09442_ net1115 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[29\] net909
+ net663 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[29\] vssd1 vssd1 vccd1
+ vccd1 _05782_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_82_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09373_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[26\] net668 _05709_ _05710_
+ _05712_ vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09231__C net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout244_A _07862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10377__C net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08324_ net990 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[30\] net951 vssd1
+ vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__and3_1
XANTENNA_wire886_X net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08255_ net2212 net2304 net1053 vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__mux2_1
XANTENNA__12365__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout411_A _03563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout509_A _06032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1153_A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08186_ net2640 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[87\] net1047 vssd1 vssd1
+ vccd1 vccd1 _03501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1320_A net1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1418_A net1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1039_X net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09980__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08431__X _04771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout780_A net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout499_X net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout878_A _04810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11709__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13513__B1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1206_X net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout666_X net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14069__B2 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09709_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[21\] net798 net731 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__a22o_1
XANTENNA__09703__A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10981_ _06905_ _07317_ _07320_ vssd1 vssd1 vccd1 vccd1 _07321_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12720_ team_01_WB.instance_to_wrap.cpu.RU0.state\[6\] team_01_WB.instance_to_wrap.cpu.RU0.state\[2\]
+ net1065 net1178 vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__o31a_1
XFILLER_0_85_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12651_ net2645 net319 net393 vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11602_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] _07818_ vssd1 vssd1
+ vccd1 vccd1 _07819_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09799__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15370_ net1295 vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12582_ net2654 net292 net401 vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__mux2_1
XANTENNA__09653__D1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14321_ net1330 vssd1 vssd1 vccd1 vccd1 _00115_ sky130_fd_sc_hd__inv_2
X_11533_ net1712 net1172 net589 net1127 vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__a22o_1
XANTENNA__12275__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14056__A _04226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17040_ clknet_leaf_144_wb_clk_i _02727_ _01023_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_11464_ _07754_ net366 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[31\] net874
+ vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__o2bb2a_1
X_14252_ net1206 vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13203_ net5 net836 net629 net2720 vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__o22a_1
X_10415_ net1133 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[27\] net982
+ vssd1 vssd1 vccd1 vccd1 _06755_ sky130_fd_sc_hd__and3_1
X_14183_ _04453_ _04454_ vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__nor2_1
XANTENNA__09420__A1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11395_ net326 _07715_ _07720_ vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10346_ net1137 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[17\] net948
+ vssd1 vssd1 vccd1 vccd1 _06686_ sky130_fd_sc_hd__and3_1
X_13134_ net1639 net845 net633 team_01_WB.instance_to_wrap.a1.ADR_I\[9\] vssd1 vssd1
+ vccd1 vccd1 _02007_ sky130_fd_sc_hd__a22o_1
X_17942_ net1457 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
X_13065_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[21\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[29\]
+ net859 vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__mux2_1
X_10277_ net1129 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[19\] net977
+ vssd1 vssd1 vccd1 vccd1 _06617_ sky130_fd_sc_hd__and3_1
XANTENNA__10318__B1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12016_ net1685 net300 net470 vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__mux2_1
Xfanout1420 net1422 vssd1 vssd1 vccd1 vccd1 net1420 sky130_fd_sc_hd__buf_2
X_17873_ clknet_leaf_127_wb_clk_i _03548_ _01813_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16824_ clknet_leaf_61_wb_clk_i _02511_ _00807_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_16755_ clknet_leaf_18_wb_clk_i _02442_ _00738_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13967_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[4\]
+ _04220_ _04223_ vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__and4_4
XANTENNA__10759__A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15706_ net1373 vssd1 vssd1 vccd1 vccd1 _01500_ sky130_fd_sc_hd__inv_2
X_12918_ net360 _03687_ net1037 vssd1 vssd1 vccd1 vccd1 _03688_ sky130_fd_sc_hd__o21ai_1
X_16686_ clknet_leaf_38_wb_clk_i _02373_ _00669_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13898_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[4\] _04141_ vssd1 vssd1 vccd1
+ vccd1 _04201_ sky130_fd_sc_hd__nand2_1
X_15637_ net1277 vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__inv_2
XANTENNA__09051__C net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12849_ net2456 net263 net381 vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10197__C net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15568_ net1274 vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08890__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17307_ clknet_leaf_71_wb_clk_i _02994_ _01290_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14519_ net1406 vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__inv_2
XANTENNA__12185__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10494__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15499_ net1395 vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__inv_2
X_08040_ net1680 net569 _04526_ team_01_WB.instance_to_wrap.cpu.f0.i\[15\] vssd1 vssd1
+ vccd1 vccd1 _03551_ sky130_fd_sc_hd__a22o_1
XANTENNA_wire581_A _06705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17238_ clknet_leaf_12_wb_clk_i _02925_ _01221_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold903 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold914 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2449 sky130_fd_sc_hd__dlygate4sd3_1
X_17169_ clknet_leaf_116_wb_clk_i _02856_ _01152_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold925 team_01_WB.instance_to_wrap.cpu.f0.num\[5\] vssd1 vssd1 vccd1 vccd1 net2460
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08899__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold936 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2471 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10021__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold947 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[43\] vssd1 vssd1 vccd1 vccd1
+ net2482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2493 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09962__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09991_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[2\] net753 net747 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06331_ sky130_fd_sc_hd__a22o_1
Xhold969 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2504 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08942_ net1026 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[6\] net931 vssd1
+ vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09175__B1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09714__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08873_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[3\] net681 _05194_ _05195_
+ _05206_ vssd1 vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_4_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1603 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net3138 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1614 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net3149 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout194_A _07634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1625 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net3160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1636 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net3171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1647 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 net3182
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout459_A _07955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10088__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09425_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[28\] net671 net660 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[28\]
+ _05762_ vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__a221o_1
XFILLER_0_137_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout626_A net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1368_A net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07978__A team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09356_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[25\] net682 _05694_
+ _05695_ vssd1 vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__a211o_1
XANTENNA__08426__X _04766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_139_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_139_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_74_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13982__B1 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08307_ net1131 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[30\] net970
+ vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09287_ net1005 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[22\] net900
+ vssd1 vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12095__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout414_X net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1156_X net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08238_ net2482 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[35\] net1054 vssd1 vssd1
+ vccd1 vccd1 _03449_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout995_A _04491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08305__C net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10548__A0 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08169_ net2860 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[104\] net1047 vssd1 vssd1
+ vccd1 vccd1 _03518_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10200_ net1142 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[8\] net963 vssd1
+ vssd1 vccd1 vccd1 _06540_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10012__A2 _04634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_152_Left_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09953__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11180_ net563 _07173_ _07510_ _07519_ vssd1 vssd1 vccd1 vccd1 _07520_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout783_X net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10131_ net372 _06467_ vssd1 vssd1 vccd1 vccd1 _06471_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_73_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08321__B net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10062_ _06399_ _06400_ _06369_ vssd1 vssd1 vccd1 vccd1 _06402_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_110_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout950_X net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09136__C net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14870_ net1246 vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_141_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13821_ net2178 net832 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[14\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_106_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16540_ clknet_leaf_6_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[6\]
+ _00523_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_13752_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[0\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[1\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[3\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__and4_2
X_10964_ _06905_ _07198_ _07300_ net531 vssd1 vssd1 vccd1 vccd1 _07304_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12703_ net2651 net262 net383 vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__mux2_1
X_16471_ clknet_leaf_140_wb_clk_i _02225_ _00454_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13683_ team_01_WB.instance_to_wrap.cpu.c0.count\[9\] _04105_ vssd1 vssd1 vccd1 vccd1
+ _04106_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08692__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10895_ net530 _07234_ vssd1 vssd1 vccd1 vccd1 _07235_ sky130_fd_sc_hd__or2_1
XANTENNA__13105__D _03728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11902__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15422_ net1350 vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__inv_2
X_12634_ net2700 net238 net391 vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13402__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15353_ net1237 vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__inv_2
X_12565_ net2247 net202 net399 vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_117_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14304_ net1330 vssd1 vssd1 vccd1 vccd1 _00098_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_117_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11516_ net1606 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[2\] team_01_WB.instance_to_wrap.cpu.DM0.next_enable
+ vssd1 vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15284_ net1379 vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__inv_2
X_12496_ net3050 net207 net409 vssd1 vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17023_ clknet_leaf_43_wb_clk_i _02710_ _01006_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14235_ net1323 vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__inv_2
X_11447_ team_01_WB.instance_to_wrap.cpu.f0.i\[3\] _07673_ net325 vssd1 vssd1 vccd1
+ vccd1 _07748_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10539__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09608__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14166_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[4\] _04188_ net1572 vssd1
+ vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__a21oi_1
X_11378_ _04475_ _07706_ vssd1 vssd1 vccd1 vccd1 _07707_ sky130_fd_sc_hd__nor2_2
XANTENNA__08512__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13117_ net1717 net846 net633 team_01_WB.instance_to_wrap.a1.ADR_I\[26\] vssd1 vssd1
+ vccd1 vccd1 _02024_ sky130_fd_sc_hd__a22o_1
X_10329_ _06646_ _06653_ _06668_ vssd1 vssd1 vccd1 vccd1 _06669_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_130_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[101\] _04254_ _04261_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[117\]
+ _04383_ vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__a221o_1
X_17925_ net1532 vssd1 vssd1 vccd1 vccd1 gpio_oeb[34] sky130_fd_sc_hd__buf_2
X_13048_ net2765 net2687 net855 vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__mux2_1
XANTENNA__09046__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1250 net1252 vssd1 vssd1 vccd1 vccd1 net1250 sky130_fd_sc_hd__buf_4
Xfanout1261 net1264 vssd1 vssd1 vccd1 vccd1 net1261 sky130_fd_sc_hd__buf_4
X_17856_ clknet_leaf_117_wb_clk_i net1821 _01796_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[126\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1272 net1273 vssd1 vssd1 vccd1 vccd1 net1272 sky130_fd_sc_hd__buf_4
Xfanout1283 net1285 vssd1 vssd1 vccd1 vccd1 net1283 sky130_fd_sc_hd__buf_4
XFILLER_0_56_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1294 net1301 vssd1 vssd1 vccd1 vccd1 net1294 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08885__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09343__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16807_ clknet_leaf_104_wb_clk_i _02494_ _00790_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_17787_ clknet_leaf_94_wb_clk_i _03463_ _01727_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[57\]
+ sky130_fd_sc_hd__dfrtp_1
X_14999_ net1213 vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16738_ clknet_leaf_75_wb_clk_i _02425_ _00721_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08407__A_N _04738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08132__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16669_ clknet_leaf_70_wb_clk_i _02356_ _00652_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12908__S net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11812__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09210_ net1085 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[17\] net939
+ vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__and3_1
XFILLER_0_57_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09141_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[14\] net651 _05458_ _05473_
+ _05479_ vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12767__A1 _07171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09072_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[12\] net655 _05385_
+ _05391_ net707 vssd1 vssd1 vccd1 vccd1 _05412_ sky130_fd_sc_hd__a2111o_1
XANTENNA_wire584_X net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08023_ team_01_WB.instance_to_wrap.cpu.f0.state\[5\] team_01_WB.instance_to_wrap.cpu.f0.state\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__nor2_1
Xhold700 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2235 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12643__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold711 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2246 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09396__B1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold722 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2257 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold733 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2279 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09935__A2 _04634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold755 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2290 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_39_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold766 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2312 sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2323 sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ net547 net534 net517 net529 vssd1 vssd1 vccd1 vccd1 _06314_ sky130_fd_sc_hd__o31a_1
Xhold799 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2334 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14141__B1 _04259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08925_ _05076_ net555 vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__or2_2
Xhold1400 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[89\] vssd1 vssd1 vccd1 vccd1
+ net2935 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1411 _03478_ vssd1 vssd1 vccd1 vccd1 net2946 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1422 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2957 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1433 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2968 sky130_fd_sc_hd__dlygate4sd3_1
X_08856_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[3\] net672 net646 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__a22o_1
Xhold1444 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2979 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08795__C net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09253__A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1455 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2990 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1466 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net3001 sky130_fd_sc_hd__dlygate4sd3_1
X_17979__1494 vssd1 vssd1 vccd1 vccd1 _17979__1494/HI net1494 sky130_fd_sc_hd__conb_1
Xhold1477 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net3012 sky130_fd_sc_hd__dlygate4sd3_1
X_08787_ net1014 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[0\] net926 vssd1
+ vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout743_A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout364_X net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1488 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net3023 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1499 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net3034 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_49_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09320__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout910_A net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09408_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[27\] net688 net656 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[27\]
+ _05747_ vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__a221o_1
X_10680_ _05901_ _06825_ _06827_ vssd1 vssd1 vccd1 vccd1 _07020_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12758__A1 _07111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09339_ net1080 net710 net594 vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_97_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09623__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_78_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_124_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12350_ net3128 net298 net430 vssd1 vssd1 vccd1 vccd1 _02645_ sky130_fd_sc_hd__mux2_1
XANTENNA__10233__A2 _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11430__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_23_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout998_X net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11301_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] _05153_ _05154_ vssd1
+ vssd1 vccd1 vccd1 _07641_ sky130_fd_sc_hd__or3_1
X_12281_ net2866 net283 net436 vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12553__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14020_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[122\] _04250_ _04268_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[74\]
+ vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__a22o_1
XANTENNA__09387__B1 _04841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11232_ _06935_ _07261_ vssd1 vssd1 vccd1 vccd1 _07572_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_112_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12930__A1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11163_ _07210_ _07255_ net516 vssd1 vssd1 vccd1 vccd1 _07503_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_36_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10114_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[6\] net820 net818 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06454_ sky130_fd_sc_hd__a22o_1
XANTENNA__14132__B1 _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11094_ _07432_ _07433_ vssd1 vssd1 vccd1 vccd1 _07434_ sky130_fd_sc_hd__nand2b_1
X_15971_ net1368 vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__inv_2
X_17710_ clknet_leaf_132_wb_clk_i _03394_ _01651_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10045_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[0\] net801 net779 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[0\]
+ _06379_ vssd1 vssd1 vccd1 vccd1 _06385_ sky130_fd_sc_hd__a221o_1
X_14922_ net1374 vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__inv_2
Xhold60 net117 vssd1 vssd1 vccd1 vccd1 net1595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[2\] vssd1 vssd1 vccd1 vccd1
+ net1606 sky130_fd_sc_hd__dlygate4sd3_1
X_17641_ clknet_leaf_0_wb_clk_i _03326_ _01582_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold82 _01994_ vssd1 vssd1 vccd1 vccd1 net1617 sky130_fd_sc_hd__dlygate4sd3_1
X_14853_ net1262 vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__inv_2
Xhold93 team_01_WB.instance_to_wrap.cpu.f0.write_data\[29\] vssd1 vssd1 vccd1 vccd1
+ net1628 sky130_fd_sc_hd__dlygate4sd3_1
X_13804_ _04158_ _01834_ _01835_ _01833_ vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__or4_1
X_17572_ clknet_leaf_87_wb_clk_i _03259_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_14784_ net1231 vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__inv_2
XANTENNA__13643__C1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11996_ net2484 net216 net468 vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__mux2_1
X_16523_ clknet_leaf_157_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[21\]
+ _00506_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13735_ _04563_ _04574_ _04503_ vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10947_ _06904_ _07281_ _07274_ _07271_ vssd1 vssd1 vccd1 vccd1 _07287_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08665__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16454_ clknet_leaf_41_wb_clk_i _02208_ _00437_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13666_ team_01_WB.instance_to_wrap.a1.WRITE_I team_01_WB.instance_to_wrap.a1.READ_I
+ vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__xnor2_1
X_10878_ _07037_ _07039_ net520 vssd1 vssd1 vccd1 vccd1 _07218_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15405_ net1263 vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__inv_2
X_12617_ net2092 net307 net398 vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_970 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16385_ clknet_leaf_97_wb_clk_i _02139_ _00368_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[108\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_115_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13597_ net988 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] _04039_ _04040_
+ vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__a22o_1
X_15336_ net1387 vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__inv_2
X_12548_ net2028 net296 net405 vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12463__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15267_ net1234 vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__inv_2
X_12479_ net2058 net281 net412 vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__mux2_1
XANTENNA_2 _03654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17006_ clknet_leaf_37_wb_clk_i _02693_ _00989_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13174__A1 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14218_ net2967 vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09917__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15198_ net1345 vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__inv_2
XANTENNA__11185__B1 _07524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12921__A1 _05528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14149_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[55\] _04262_ _04266_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[23\]
+ _04152_ vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__a221o_1
Xfanout509 _06032_ vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14123__B1 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08710_ net1102 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[5\] net932 vssd1
+ vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__and3_1
XANTENNA__11807__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17908_ net1519 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
X_09690_ _06019_ _06024_ _06029_ vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__or3_2
Xfanout1080 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[24\] vssd1 vssd1 vccd1 vccd1
+ net1080 sky130_fd_sc_hd__clkbuf_8
X_08641_ net1021 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[10\] net927 vssd1
+ vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__and3_1
Xfanout1091 net1096 vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__buf_1
XFILLER_0_20_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17839_ clknet_leaf_97_wb_clk_i _03515_ _01779_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[109\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__09504__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08572_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[19\] net658 _04909_
+ _04910_ _04911_ vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_117_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08656__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_112_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12638__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11660__A1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10463__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08417__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout324_A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1066_A net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10215__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09124_ net1104 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[14\] net889
+ vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__and3_1
XANTENNA_wire966_X net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09055_ net1110 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[12\] net902
+ vssd1 vssd1 vccd1 vccd1 _05395_ sky130_fd_sc_hd__and3_1
XFILLER_0_130_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12373__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1233_A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13165__A1 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09369__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08006_ team_01_WB.instance_to_wrap.cpu.f0.state\[2\] vssd1 vssd1 vccd1 vccd1 _04503_
+ sky130_fd_sc_hd__inv_2
Xhold530 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2065 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11497__B _07756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout693_A _04771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold541 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2076 sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2087 sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 team_01_WB.instance_to_wrap.cpu.c0.count\[14\] vssd1 vssd1 vccd1 vccd1 net2098
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[6\] vssd1 vssd1 vccd1 vccd1
+ net2109 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1021_X net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1400_A net1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold585 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2131 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07991__A team_01_WB.instance_to_wrap.cpu.f0.i\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14114__B1 _04236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09957_ net1155 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[3\] net969 vssd1
+ vssd1 vccd1 vccd1 _06297_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout481_X net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout860_A net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout958_A net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08908_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[2\] net695 _05225_ _05241_
+ _05242_ vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__a2111o_1
X_09888_ net1153 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[5\] net985 vssd1
+ vssd1 vccd1 vccd1 _06228_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_151_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold1230 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[38\] vssd1 vssd1 vccd1 vccd1
+ net2765 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1241 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1252 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2787 sky130_fd_sc_hd__dlygate4sd3_1
X_08839_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[1\] net687 _05161_ _05167_
+ net706 vssd1 vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__a2111o_1
Xhold1263 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2798 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1274 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2809 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout746_X net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1285 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2820 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1296 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2831 sky130_fd_sc_hd__dlygate4sd3_1
X_11850_ net2435 net301 net488 vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_154_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_154_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_131_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10801_ net522 _06972_ _07140_ vssd1 vssd1 vccd1 vccd1 _07141_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_67_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12548__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11781_ net2090 net280 net497 vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout913_X net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13640__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13520_ _03851_ _03943_ _03850_ vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_64_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10732_ _05781_ _05898_ vssd1 vssd1 vccd1 vccd1 _07072_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_24_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08327__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13451_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] _05381_ _05419_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\]
+ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10663_ _07001_ _07002_ net541 vssd1 vssd1 vccd1 vccd1 _07003_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12402_ net2571 net269 net419 vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__mux2_1
X_16170_ clknet_leaf_3_wb_clk_i _00012_ _00158_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_153_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10594_ net553 _06902_ vssd1 vssd1 vccd1 vccd1 _06934_ sky130_fd_sc_hd__nor2_2
X_13382_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] _05803_ vssd1 vssd1
+ vccd1 vccd1 _03843_ sky130_fd_sc_hd__nand2_1
XANTENNA__09072__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15121_ net1422 vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__inv_2
XANTENNA__10757__A3 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08280__A0 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12333_ net2599 net203 net427 vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__mux2_1
XANTENNA__12283__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15052_ net1265 vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09158__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12264_ net2833 net247 net437 vssd1 vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14003_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[25\] _04243_ _04268_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[73\]
+ vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__a22o_1
XANTENNA__12903__A1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11706__A2 _07531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16052__Q team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11215_ _06750_ _06817_ _06822_ vssd1 vssd1 vccd1 vccd1 _07555_ sky130_fd_sc_hd__a21oi_2
XANTENNA__10914__A0 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12195_ net2453 net210 net443 vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__mux2_1
XANTENNA__14105__B1 _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09780__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__buf_2
X_11146_ _06920_ _07241_ _07275_ _07238_ vssd1 vssd1 vccd1 vccd1 _07486_ sky130_fd_sc_hd__o211a_1
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 ADR_O[27] sky130_fd_sc_hd__buf_2
XANTENNA__11627__S net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11077_ net505 _04919_ vssd1 vssd1 vccd1 vccd1 _07417_ sky130_fd_sc_hd__and2b_1
X_15954_ net1363 vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_129_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10028_ net561 net552 net535 vssd1 vssd1 vccd1 vccd1 _06368_ sky130_fd_sc_hd__o21ai_1
X_14905_ net1238 vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__inv_2
X_15885_ net1415 vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17624_ clknet_leaf_5_wb_clk_i _03309_ _01565_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\]
+ sky130_fd_sc_hd__dfrtp_2
X_14836_ net1399 vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17555_ clknet_leaf_16_wb_clk_i _03242_ _01538_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_14767_ net1385 vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__inv_2
XANTENNA__12458__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11979_ net2163 net284 net473 vssd1 vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__mux2_1
XANTENNA__14239__A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16506_ clknet_leaf_6_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[4\]
+ _00489_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13718_ _04105_ _04128_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[8\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_156_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17486_ clknet_leaf_38_wb_clk_i _03173_ _01469_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14698_ net1210 vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16437_ clknet_leaf_49_wb_clk_i _02191_ _00420_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13649_ net727 _07507_ net988 vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16368_ clknet_leaf_97_wb_clk_i net1543 _00351_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[91\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15319_ net1221 vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__inv_2
XANTENNA__12193__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16299_ clknet_leaf_125_wb_clk_i net2621 _00282_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_17978__1493 vssd1 vssd1 vccd1 vccd1 _17978__1493/HI net1493 sky130_fd_sc_hd__conb_1
XANTENNA__08810__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_779 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13552__D1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout306 _07935_ vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout317 net320 vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__buf_2
X_09811_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[14\] net773 net737 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06151_ sky130_fd_sc_hd__a22o_1
XANTENNA__11173__A3 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09771__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout328 _07070_ vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__clkbuf_4
Xfanout339 _06590_ vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__clkbuf_4
X_09742_ net1145 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[20\] net964
+ vssd1 vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__and3_1
XANTENNA__09523__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09673_ net1135 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[22\] net945
+ vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__and3_1
XANTENNA__08877__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08624_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[11\] net676 net661 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[11\]
+ _04954_ vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__a221o_1
XANTENNA__13607__C1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13083__A0 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09531__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08555_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[19\] net654 net652 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[19\]
+ _04894_ vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__a221o_1
XANTENNA__08629__A2 _04968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout441_A _07962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12368__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1183_A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08418__Y _04758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13622__A2 _07531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11633__A1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10436__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08486_ net1082 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[23\] net940
+ vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__and3_1
XFILLER_0_108_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12892__A _05678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1350_A net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout706_A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout327_X net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1069_X net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09107_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[13\] net646 _05428_
+ _05435_ _05437_ vssd1 vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_131_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11301__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09038_ _05264_ _05265_ _05302_ _05377_ vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__nor4b_2
XFILLER_0_131_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout696_X net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11020__B net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15708__A net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold360 team_01_WB.instance_to_wrap.a1.ADR_I\[19\] vssd1 vssd1 vccd1 vccd1 net1895
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 team_01_WB.instance_to_wrap.cpu.f0.i\[27\] vssd1 vssd1 vccd1 vccd1 net1906
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12897__B1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold382 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1917 sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1928 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ _06974_ _06975_ _06883_ vssd1 vssd1 vccd1 vccd1 _07340_ sky130_fd_sc_hd__o21ba_1
XANTENNA__09706__A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout840 net841 vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__buf_2
Xfanout851 _03731_ vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__buf_4
XFILLER_0_99_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout862 net867 vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__clkbuf_2
Xfanout873 _00017_ vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__clkbuf_4
Xfanout884 net885 vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__buf_4
XANTENNA__09514__B1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout895 _04796_ vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__buf_4
X_12951_ net1689 net870 net357 _03710_ vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__a22o_1
XANTENNA__10959__A2_N net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10124__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1060 _02097_ vssd1 vssd1 vccd1 vccd1 net2595 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08868__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1071 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2606 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11902_ net1784 net201 net479 vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__mux2_1
X_15670_ net1247 vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__inv_2
XANTENNA__11872__A1 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1082 _03454_ vssd1 vssd1 vccd1 vccd1 net2617 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1093 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[23\] vssd1 vssd1 vccd1 vccd1
+ net2628 sky130_fd_sc_hd__dlygate4sd3_1
X_12882_ net1835 net869 net356 _03662_ vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__a22o_1
XANTENNA__08983__C net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14621_ net1323 vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__inv_2
X_11833_ net3146 net207 net489 vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12278__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13613__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17340_ clknet_leaf_58_wb_clk_i _03027_ _01323_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_14552_ net1352 vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__inv_2
XANTENNA__10427__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12821__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11764_ net2924 net247 net496 vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_155_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13503_ net987 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] _03961_ _03962_
+ vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__a22o_1
XANTENNA__16047__Q team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10715_ net553 _06928_ vssd1 vssd1 vccd1 vccd1 _07055_ sky130_fd_sc_hd__nand2_1
X_17271_ clknet_leaf_14_wb_clk_i _02958_ _01254_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_14483_ net1417 vssd1 vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__inv_2
X_11695_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[12\] net714 vssd1 vssd1 vccd1
+ vccd1 _07893_ sky130_fd_sc_hd__or2_1
XANTENNA__11910__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16222_ clknet_leaf_139_wb_clk_i net1580 _00210_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__dfrtp_1
XANTENNA__13377__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13434_ _03893_ _03894_ vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10646_ net509 net508 net543 vssd1 vssd1 vccd1 vccd1 _06986_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11388__B1 _07699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16153_ clknet_leaf_131_wb_clk_i _01916_ _00141_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13410__B _05220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13365_ net586 _07683_ _03834_ net565 _04485_ vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_51_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10577_ _04741_ _04744_ vssd1 vssd1 vccd1 vccd1 _06917_ sky130_fd_sc_hd__or2_2
XFILLER_0_2_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15104_ net1234 vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__inv_2
X_12316_ net2286 net278 net432 vssd1 vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__mux2_1
X_16084_ clknet_leaf_131_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[6\]
+ _00072_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[6\] sky130_fd_sc_hd__dfrtp_1
X_13296_ _07650_ _03779_ _03781_ net825 net1540 vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__o32a_1
XFILLER_0_146_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15035_ net1250 vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__inv_2
X_12247_ net2165 net250 net442 vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__mux2_1
XANTENNA__12741__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12888__B1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_39_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12178_ net2736 net225 net447 vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__mux2_1
X_11129_ _07466_ _07468_ net554 vssd1 vssd1 vccd1 vccd1 _07469_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16986_ clknet_leaf_78_wb_clk_i _02673_ _00969_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_127_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09054__C net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15937_ net1402 vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15868_ net1202 vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__inv_2
XANTENNA__08666__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08893__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17607_ clknet_leaf_86_wb_clk_i _03294_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_14819_ net1250 vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__inv_2
XANTENNA__12188__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15799_ net1230 vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08340_ net1155 net953 vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__and2_2
X_17538_ clknet_leaf_56_wb_clk_i _03225_ _01521_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12812__B1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08271_ net2224 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[2\] net1053 vssd1 vssd1
+ vccd1 vccd1 _03416_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17469_ clknet_leaf_69_wb_clk_i _03156_ _01452_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11091__A2 _06882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13368__A1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11820__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11121__A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10051__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12651__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12879__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08701__Y _05041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1029_A net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09744__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout391_A net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout489_A _07947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07986_ team_01_WB.instance_to_wrap.cpu.f0.i\[9\] vssd1 vssd1 vccd1 vccd1 _04484_
+ sky130_fd_sc_hd__inv_2
XANTENNA__14096__A2 _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09725_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] net626 _06063_ _06064_
+ vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_87_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout656_A _04815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1398_A net1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09656_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] net625 _05994_ _05995_
+ vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_2_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08607_ _04944_ _04945_ net597 vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__mux2_2
XANTENNA__12098__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout823_A net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09587_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[25\] net735 _05908_ _05910_
+ _05914_ vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout444_X net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08538_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[18\] net690 _04849_ _04863_
+ net705 vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12803__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09275__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11015__B net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout611_X net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12826__S net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08469_ net1002 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[23\] net901
+ vssd1 vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11730__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10500_ net1130 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[31\] net972
+ vssd1 vssd1 vccd1 vccd1 _06840_ sky130_fd_sc_hd__and3b_1
XFILLER_0_93_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09027__A2 _04771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11480_ net366 _07767_ net2628 net874 vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_150_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14020__A2 _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_150_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10431_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[27\] net745 net734 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06771_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09983__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13150_ net126 net847 net839 net1609 vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_59_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10362_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[17\] net816 net794 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _06702_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_59_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout980_X net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09139__C net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12101_ net1918 net200 net455 vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__mux2_1
XANTENNA__12561__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10293_ _06627_ _06628_ _06632_ vssd1 vssd1 vccd1 vccd1 _06633_ sky130_fd_sc_hd__or3_1
X_13081_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[13\]
+ net860 vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08978__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12032_ net3059 net208 net465 vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__mux2_1
XANTENNA__13531__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold190 team_01_WB.instance_to_wrap.a1.ADR_I\[15\] vssd1 vssd1 vccd1 vccd1 net1725
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11685__B net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08340__A net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16840_ clknet_leaf_62_wb_clk_i _02527_ _00823_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout670 _04800_ vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__buf_8
Xfanout681 _04787_ vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__buf_4
XANTENNA__09723__X _06063_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16771_ clknet_leaf_25_wb_clk_i _02458_ _00754_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout692 net693 vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13295__B1 _04621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13983_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[112\] _04261_ _04262_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[48\]
+ _04274_ vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__a221o_1
XANTENNA__11905__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15722_ net1283 vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__inv_2
X_12934_ _05415_ _07757_ _03694_ vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_137_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10588__Y _06928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17977__1492 vssd1 vssd1 vccd1 vccd1 _17977__1492/HI net1492 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_122_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09171__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15653_ net1262 vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__inv_2
X_12865_ net2088 net288 net382 vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__mux2_1
XANTENNA__13405__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09602__C net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13598__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14604_ net1329 vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__inv_2
X_11816_ net1833 net278 net492 vssd1 vssd1 vccd1 vccd1 _03158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15584_ net1230 vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__inv_2
X_12796_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] net1060 net363 _03625_
+ vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__a22o_1
XANTENNA__09266__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17323_ clknet_leaf_9_wb_clk_i _03010_ _01306_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14535_ net1406 vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__inv_2
XANTENNA__10805__C1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11747_ net2149 net307 net500 vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17254_ clknet_leaf_83_wb_clk_i _02941_ _01237_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14466_ net1357 vssd1 vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__inv_2
X_11678_ _07878_ _07879_ net612 vssd1 vssd1 vccd1 vccd1 _07880_ sky130_fd_sc_hd__mux2_4
XANTENNA__14011__A2 _04246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16205_ clknet_leaf_140_wb_clk_i _01965_ _00193_ vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__dfrtp_2
XFILLER_0_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13417_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] _05112_ vssd1 vssd1 vccd1
+ vccd1 _03878_ sky130_fd_sc_hd__or2_1
X_17185_ clknet_leaf_52_wb_clk_i _02872_ _01168_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10629_ net537 _06968_ vssd1 vssd1 vccd1 vccd1 _06969_ sky130_fd_sc_hd__nand2_2
XFILLER_0_107_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14397_ net1189 vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10033__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16136_ clknet_leaf_158_wb_clk_i _00010_ _00124_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.curr_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09974__B1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13348_ net565 _07680_ _03819_ _03821_ vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_47_Left_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09049__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12471__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16067_ clknet_leaf_157_wb_clk_i _01860_ _00055_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10780__A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13279_ team_01_WB.instance_to_wrap.cpu.f0.i\[26\] _03753_ vssd1 vssd1 vccd1 vccd1
+ _03768_ sky130_fd_sc_hd__nand2_1
XANTENNA__14252__A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12324__X _07965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08888__C net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15018_ net1283 vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__inv_2
XANTENNA__13522__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11595__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14078__A2 _04236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16969_ clknet_leaf_40_wb_clk_i _02656_ _00952_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11815__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09510_ net1150 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[29\] net959
+ vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_56_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08701__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09441_ _05779_ _05780_ net598 vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_82_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13589__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09372_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[26\] net657 net655 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[26\]
+ _05711_ vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__a221o_1
XANTENNA__09257__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08323_ net991 net951 vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__and2_1
XANTENNA__12646__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout237_A net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08254_ net2587 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[19\] net1055 vssd1 vssd1
+ vccd1 vccd1 _03433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14002__A2 _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12013__A1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13210__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08185_ net2956 net2876 net1047 vssd1 vssd1 vccd1 vccd1 _03502_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_65_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout404_A net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1146_A net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_924 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12381__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13513__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09717__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08798__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09256__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout394_X net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout773_A net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1101_X net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14069__A2 _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07969_ team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1 _04467_
+ sky130_fd_sc_hd__inv_2
XANTENNA_fanout561_X net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout940_A _04759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_74_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11725__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout659_X net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09708_ net1148 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[21\] net946
+ vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_143_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10980_ net531 _07182_ _07319_ net375 vssd1 vssd1 vccd1 vccd1 _07320_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09639_ net1135 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[23\] net954
+ vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__and3_1
XANTENNA__08319__B net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12650_ net2461 net305 net392 vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__mux2_1
XANTENNA__09248__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11601_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\]
+ _07817_ vssd1 vssd1 vccd1 vccd1 _07818_ sky130_fd_sc_hd__and3_1
XFILLER_0_93_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12581_ net2525 net299 net402 vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__mux2_1
XANTENNA__12556__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14320_ net1348 vssd1 vssd1 vccd1 vccd1 _00114_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11532_ net1740 net1171 net589 net1124 vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_83_Left_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14056__B _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14251_ net1206 vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__inv_2
XANTENNA__13201__B1 _03738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11463_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[15\] _07755_ _07758_ vssd1 vssd1
+ vccd1 vccd1 _07759_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_78_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire378 team_01_WB.instance_to_wrap.cpu.RU0.next_write_i vssd1 vssd1 vccd1 vccd1
+ net378 sky130_fd_sc_hd__clkbuf_2
X_13202_ net6 net835 net628 net1708 vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_78_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10015__B1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10414_ net1132 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[27\] net975
+ vssd1 vssd1 vccd1 vccd1 _06754_ sky130_fd_sc_hd__and3_1
X_14182_ net2103 _04452_ net1183 vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11394_ net1068 _07668_ _07714_ team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1
+ vssd1 vccd1 vccd1 _07720_ sky130_fd_sc_hd__a31o_1
XFILLER_0_61_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13133_ net76 net844 net632 net1630 vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__a22o_1
X_10345_ net1137 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[17\] net958
+ vssd1 vssd1 vccd1 vccd1 _06685_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_115_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09166__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17941_ net1456 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
XFILLER_0_40_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13064_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[22\] net2846 net853 vssd1 vssd1
+ vccd1 vccd1 _02061_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10276_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[19\] net745 _06613_ _06614_
+ _06615_ vssd1 vssd1 vccd1 vccd1 _06616_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10318__A1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16060__Q team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12015_ net1860 net280 net470 vssd1 vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__mux2_1
Xfanout1410 net1414 vssd1 vssd1 vccd1 vccd1 net1410 sky130_fd_sc_hd__buf_4
Xfanout1421 net1422 vssd1 vssd1 vccd1 vccd1 net1421 sky130_fd_sc_hd__buf_4
X_17872_ clknet_leaf_115_wb_clk_i _03547_ _01812_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_16823_ clknet_leaf_11_wb_clk_i _02510_ _00806_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16754_ clknet_leaf_143_wb_clk_i _02441_ _00737_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13966_ _04238_ _04257_ vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_17_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12917_ _05564_ net577 vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__nor2_1
X_15705_ net1240 vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__inv_2
X_16685_ clknet_leaf_108_wb_clk_i _02372_ _00668_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13897_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[4\] _04141_ vssd1 vssd1 vccd1
+ vccd1 _04200_ sky130_fd_sc_hd__or2_1
XFILLER_0_152_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12848_ net3091 net265 net382 vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__mux2_1
X_15636_ net1399 vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__inv_2
XANTENNA__09239__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15567_ net1299 vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12466__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13862__A_N net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12779_ net1545 net638 net606 _03614_ vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_79 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08998__A1 _05337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17306_ clknet_leaf_78_wb_clk_i _02993_ _01289_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14518_ net1354 vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__inv_2
X_15498_ net1377 vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14449_ net1225 vssd1 vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__inv_2
X_17237_ clknet_leaf_109_wb_clk_i _02924_ _01220_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17168_ clknet_leaf_146_wb_clk_i _02855_ _01151_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold904 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2439 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17464__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold915 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2450 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09411__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold926 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold937 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2472 sky130_fd_sc_hd__dlygate4sd3_1
X_16119_ clknet_leaf_134_wb_clk_i _01894_ _00107_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_29_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold948 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2483 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09990_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[2\] net805 net750 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06330_ sky130_fd_sc_hd__a22o_1
Xhold959 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2494 sky130_fd_sc_hd__dlygate4sd3_1
X_17099_ clknet_leaf_8_wb_clk_i _02786_ _01082_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_08941_ net1028 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[6\] net920 vssd1
+ vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__and3_1
XANTENNA__09507__C net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09175__A1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15806__A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_wb_clk_i_A wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08872_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[3\] _04806_ _05198_
+ _05200_ _05202_ vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_32_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1604 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[15\] vssd1 vssd1 vccd1 vccd1
+ net3139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1615 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net3150 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1626 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net3161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1637 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 net3172
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1648 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1 net3183
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout187_A _07639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09478__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1096_A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09424_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[28\] net688 net646 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[28\]
+ _05763_ vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09355_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[25\] net669 net651 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__a22o_1
XANTENNA__12376__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout521_A _05260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10245__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08306_ net1155 net970 vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__and2_2
XANTENNA_clkbuf_leaf_68_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09286_ net1004 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[22\] net888 vssd1
+ vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08237_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[44\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[36\]
+ net1050 vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1430_A net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout407_X net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07994__A team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08168_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[113\] net2403 net1056 vssd1 vssd1
+ vccd1 vccd1 _03519_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout890_A _04799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10548__A1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09402__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_108_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_108_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_132_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout988_A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17976__1491 vssd1 vssd1 vccd1 vccd1 _17976__1491/HI net1491 sky130_fd_sc_hd__conb_1
XANTENNA__08610__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08099_ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[0\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10130_ _06438_ _06440_ vssd1 vssd1 vccd1 vccd1 _06470_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_73_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout776_X net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10061_ _06369_ _06400_ vssd1 vssd1 vccd1 vccd1 _06401_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_110_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout943_X net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17704__Q team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_138_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13820_ net1708 net832 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[13\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_98_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13751_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[0\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[1\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[2\] vssd1 vssd1 vccd1 vccd1 _04140_
+ sky130_fd_sc_hd__nand3_1
XFILLER_0_97_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10963_ net539 _06940_ _06942_ _07302_ vssd1 vssd1 vccd1 vccd1 _07303_ sky130_fd_sc_hd__o31a_1
XANTENNA__13670__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12702_ net2491 net268 net383 vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__mux2_1
X_16470_ clknet_leaf_141_wb_clk_i _02224_ _00453_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13682_ team_01_WB.instance_to_wrap.cpu.c0.count\[8\] team_01_WB.instance_to_wrap.cpu.c0.count\[7\]
+ _04103_ vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__and3_1
X_10894_ _07137_ _07181_ net514 vssd1 vssd1 vccd1 vccd1 _07234_ sky130_fd_sc_hd__mux2_1
X_15421_ net1315 vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__inv_2
X_12633_ net2624 net269 net391 vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__mux2_1
XANTENNA__12286__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14067__A net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10236__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15352_ net1215 vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12564_ net2707 net205 net399 vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__mux2_1
XANTENNA__13402__C net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09641__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14303_ net1328 vssd1 vssd1 vccd1 vccd1 _00097_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16055__Q team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11515_ net1624 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[3\] net877 vssd1 vssd1
+ vccd1 vccd1 _03334_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15283_ net1383 vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12495_ net2323 net247 net409 vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__mux2_1
X_17022_ clknet_leaf_84_wb_clk_i _02709_ _01005_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09929__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14234_ net1323 vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__inv_2
XANTENNA_input72_X net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11446_ team_01_WB.instance_to_wrap.cpu.f0.i\[4\] _07674_ _07747_ vssd1 vssd1 vccd1
+ vccd1 _03367_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_145_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14165_ _04195_ _04443_ net1426 vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08601__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11377_ team_01_WB.instance_to_wrap.cpu.f0.i\[18\] _07705_ vssd1 vssd1 vccd1 vccd1
+ _07706_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13116_ net1596 net844 net631 team_01_WB.instance_to_wrap.a1.ADR_I\[27\] vssd1 vssd1
+ vccd1 vccd1 _02025_ sky130_fd_sc_hd__a22o_1
X_10328_ _06657_ _06659_ _06663_ _06667_ vssd1 vssd1 vccd1 vccd1 _06668_ sky130_fd_sc_hd__or4_1
X_14096_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[69\] _04233_ _04253_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17924_ net1531 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
X_13047_ net2602 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[47\] net857 vssd1 vssd1
+ vccd1 vccd1 _02078_ sky130_fd_sc_hd__mux2_1
X_10259_ _06193_ _06218_ _06192_ vssd1 vssd1 vccd1 vccd1 _06599_ sky130_fd_sc_hd__a21o_1
Xfanout1240 net1241 vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__buf_4
XFILLER_0_56_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1251 net1252 vssd1 vssd1 vccd1 vccd1 net1251 sky130_fd_sc_hd__buf_2
Xfanout1262 net1264 vssd1 vssd1 vccd1 vccd1 net1262 sky130_fd_sc_hd__buf_4
X_17855_ clknet_leaf_98_wb_clk_i _03531_ _01795_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[125\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout1273 net1302 vssd1 vssd1 vccd1 vccd1 net1273 sky130_fd_sc_hd__buf_2
Xfanout1284 net1285 vssd1 vssd1 vccd1 vccd1 net1284 sky130_fd_sc_hd__buf_2
Xfanout1295 net1301 vssd1 vssd1 vccd1 vccd1 net1295 sky130_fd_sc_hd__buf_4
X_16806_ clknet_leaf_72_wb_clk_i _02493_ _00789_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_17786_ clknet_leaf_123_wb_clk_i _03462_ _01726_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[56\]
+ sky130_fd_sc_hd__dfrtp_1
X_14998_ net1256 vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16737_ clknet_leaf_55_wb_clk_i _02424_ _00720_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09062__C net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13949_ _04218_ _04229_ vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__nor2_4
XANTENNA_clkbuf_leaf_102_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16668_ clknet_leaf_57_wb_clk_i _02355_ _00651_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12196__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15619_ net1252 vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16599_ clknet_leaf_15_wb_clk_i _02286_ _00582_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09140_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[14\] net697 _05461_
+ _05462_ _05468_ vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_6_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_115_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09071_ _05407_ _05408_ _05409_ _05410_ vssd1 vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__or4_2
XFILLER_0_114_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08022_ _04505_ _04516_ vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__or2_2
XFILLER_0_47_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold701 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[91\] vssd1 vssd1 vccd1 vccd1
+ net2236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold712 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2247 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11727__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold723 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2258 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13192__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold734 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2280 sky130_fd_sc_hd__dlygate4sd3_1
Xhold756 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2291 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold767 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2313 sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] net626 _06311_ _06312_
+ vssd1 vssd1 vccd1 vccd1 _06313_ sky130_fd_sc_hd__a22o_4
Xhold789 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2324 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10950__A1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08924_ net547 net534 net529 net517 vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_90_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1011_A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1109_A net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1401 team_01_WB.instance_to_wrap.cpu.f0.num\[25\] vssd1 vssd1 vccd1 vccd1 net2936
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_141_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09534__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08855_ net1024 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[3\] net919 vssd1
+ vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__and3_1
Xhold1412 team_01_WB.instance_to_wrap.cpu.f0.num\[23\] vssd1 vssd1 vccd1 vccd1 net2947
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout471_A _07952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1423 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[27\] vssd1 vssd1 vccd1 vccd1
+ net2958 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1434 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2969 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1445 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2980 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout569_A net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1456 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2991 sky130_fd_sc_hd__dlygate4sd3_1
X_08786_ net1094 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[0\] net887 vssd1
+ vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__and3_1
Xhold1467 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net3002 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1478 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net3013 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1489 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net3024 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1380_A net1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09320__A1 net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1099_X net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10466__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07989__A team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09871__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09407_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[27\] net661 net654 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout903_A _04788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09700__C net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09338_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[24\] net703 _05672_ _05677_
+ vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__o22a_4
XFILLER_0_146_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10769__A1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09623__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12834__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09269_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[20\] net672 net655 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[20\]
+ _05608_ vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__a221o_1
XFILLER_0_105_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11300_ _05153_ _05154_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] vssd1
+ vssd1 vccd1 vccd1 _07640_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_134_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12280_ net2145 net250 net437 vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout893_X net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09387__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11231_ _07569_ _07570_ vssd1 vssd1 vccd1 vccd1 _07571_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_112_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08332__B net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11162_ _07382_ _07501_ _07042_ _07101_ vssd1 vssd1 vccd1 vccd1 _07502_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_140_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10113_ _06449_ _06450_ _06451_ _06452_ vssd1 vssd1 vccd1 vccd1 _06453_ sky130_fd_sc_hd__or4_1
XANTENNA__14132__B2 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11093_ net534 _06366_ vssd1 vssd1 vccd1 vccd1 _07433_ sky130_fd_sc_hd__nand2_1
X_15970_ net1363 vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__inv_2
XANTENNA__08986__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input32_A DAT_I[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09444__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14921_ net1288 vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__inv_2
X_10044_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[0\] net752 _06373_ _06383_
+ vssd1 vssd1 vccd1 vccd1 _06384_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_76_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold50 team_01_WB.instance_to_wrap.a1.ADR_I\[24\] vssd1 vssd1 vccd1 vccd1 net1585
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 net94 vssd1 vssd1 vccd1 vccd1 net1596 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08362__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17640_ clknet_leaf_0_wb_clk_i _03325_ _01581_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold72 net78 vssd1 vssd1 vccd1 vccd1 net1607 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 net122 vssd1 vssd1 vccd1 vccd1 net1618 sky130_fd_sc_hd__dlygate4sd3_1
X_14852_ net1218 vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold94 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[30\] vssd1 vssd1 vccd1 vccd1
+ net1629 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13803_ _04159_ _04181_ _04182_ _04154_ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__a22o_1
X_17571_ clknet_leaf_87_wb_clk_i _03258_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_14783_ net1317 vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__inv_2
X_11995_ net2000 net218 net468 vssd1 vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__mux2_1
XANTENNA_output119_A net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10457__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11913__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16522_ clknet_leaf_0_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[20\]
+ _00505_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13734_ team_01_WB.instance_to_wrap.cpu.f0.state\[5\] _04516_ _04524_ _04134_ vssd1
+ vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_11_Left_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10946_ _07284_ _07285_ net521 vssd1 vssd1 vccd1 vccd1 _07286_ sky130_fd_sc_hd__mux2_1
XANTENNA__09862__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16453_ clknet_leaf_62_wb_clk_i _02207_ _00436_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13665_ net989 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] _04095_ _04096_
+ vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10877_ net558 _07216_ vssd1 vssd1 vccd1 vccd1 _07217_ sky130_fd_sc_hd__or2_1
XFILLER_0_156_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10209__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11214__A _07171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15404_ net1257 vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__inv_2
X_12616_ net2139 net311 net398 vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__mux2_1
XANTENNA__12749__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16384_ clknet_leaf_95_wb_clk_i _02138_ _00367_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[107\]
+ sky130_fd_sc_hd__dfrtp_1
X_13596_ net721 _07188_ net1075 vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09614__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_982 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15335_ net1387 vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12547_ net3154 net276 net406 vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__mux2_1
XANTENNA__12744__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15266_ net1318 vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__inv_2
X_12478_ net3064 net250 net414 vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__mux2_1
XANTENNA_3 _03654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08523__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14217_ net3072 vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__clkbuf_1
X_17005_ clknet_leaf_68_wb_clk_i _02692_ _00988_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11429_ net324 _07738_ _07739_ vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_20_Left_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15197_ net1313 vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11185__B2 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10491__C net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12921__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14148_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[15\] _04226_ _04260_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[63\]
+ _04432_ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__a221o_1
XANTENNA__08810__X _05150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09057__C net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14079_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[28\] _04243_ _04245_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[84\]
+ _04366_ vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__a221o_1
XANTENNA__14260__A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08896__C net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17907_ net1518 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
XFILLER_0_83_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1070 team_01_WB.instance_to_wrap.cpu.f0.i\[8\] vssd1 vssd1 vccd1 vccd1 net1070
+ sky130_fd_sc_hd__buf_2
X_08640_ net1100 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[10\] net893
+ vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__and3_1
Xfanout1081 net1089 vssd1 vssd1 vccd1 vccd1 net1081 sky130_fd_sc_hd__clkbuf_2
Xfanout1092 net1093 vssd1 vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__clkbuf_2
X_17838_ clknet_leaf_119_wb_clk_i _03514_ _01778_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[108\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_83_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08571_ net999 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[19\] net906 vssd1
+ vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__and3_1
XANTENNA__12437__A1 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13634__B1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17769_ clknet_leaf_121_wb_clk_i _03445_ _01709_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11823__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17975__1490 vssd1 vssd1 vccd1 vccd1 _17975__1490/HI net1490 sky130_fd_sc_hd__conb_1
XFILLER_0_77_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08417__B net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09123_ net1110 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[14\] net931
+ vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09054_ net1027 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[12\] net899 vssd1
+ vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__and3_1
XANTENNA__09529__A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08005_ team_01_WB.instance_to_wrap.cpu.c0.count\[16\] vssd1 vssd1 vccd1 vccd1 _04502_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_41_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13165__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold520 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 net2055
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2066 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08152__B net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1226_A net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold542 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 net2077
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold553 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2088 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12912__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold564 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2099 sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2110 sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2121 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold597 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 net2132
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout686_A _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08592__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09956_ net1154 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[3\] net966 vssd1
+ vssd1 vccd1 vccd1 _06296_ sky130_fd_sc_hd__and3_1
XANTENNA__08579__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1014_X net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08907_ net1026 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[2\] net880 vssd1
+ vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__and3_1
X_09887_ net998 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[5\] net969 vssd1
+ vssd1 vccd1 vccd1 _06227_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout474_X net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout853_A net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1220 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2755 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1231 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2766 sky130_fd_sc_hd__dlygate4sd3_1
X_08838_ _05175_ _05176_ _05177_ vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__or3_1
Xhold1242 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2777 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1253 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2788 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_142_Right_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1264 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[81\] vssd1 vssd1 vccd1 vccd1
+ net2799 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10151__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1275 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2810 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1286 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2821 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11018__B _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08769_ _05105_ _05106_ _05107_ _05108_ vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__or4_1
Xhold1297 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[56\] vssd1 vssd1 vccd1 vccd1
+ net2832 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1383_X net1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout739_X net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10439__B1 _06777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10800_ net524 _07139_ vssd1 vssd1 vccd1 vccd1 _07140_ sky130_fd_sc_hd__nand2_1
X_11780_ net2270 net251 net497 vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_3__f_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09844__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10731_ net553 _07069_ vssd1 vssd1 vccd1 vccd1 _07071_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_64_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout906_X net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08327__B net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13450_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] _04946_ _03910_ vssd1
+ vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__o21a_1
X_10662_ _06526_ net339 net546 vssd1 vssd1 vccd1 vccd1 _07002_ sky130_fd_sc_hd__mux2_1
XANTENNA__14050__B1 _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_123_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_123_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12401_ net2496 net243 net421 vssd1 vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__mux2_1
X_13381_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] _05803_ vssd1 vssd1
+ vccd1 vccd1 _03842_ sky130_fd_sc_hd__or2_1
XANTENNA__12564__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10593_ net557 _06930_ _06931_ _06932_ vssd1 vssd1 vccd1 vccd1 _06933_ sky130_fd_sc_hd__o22ai_1
XANTENNA__10873__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15120_ net1271 vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_11_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12332_ net2122 net272 net429 vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08343__A net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15051_ net1397 vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__inv_2
X_12263_ net3140 net213 net435 vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14002_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[49\] _04262_ _04267_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11214_ _07171_ _07207_ _07251_ _07542_ vssd1 vssd1 vccd1 vccd1 _07554_ sky130_fd_sc_hd__or4_1
XANTENNA__08032__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12194_ net3108 net214 net445 vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__mux2_1
XANTENNA__10914__A1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11908__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11145_ _05263_ _07484_ vssd1 vssd1 vccd1 vccd1 _07485_ sky130_fd_sc_hd__or2_1
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__buf_2
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__buf_2
X_11076_ _04884_ _06672_ _07127_ vssd1 vssd1 vccd1 vccd1 _07416_ sky130_fd_sc_hd__and3_1
XANTENNA__13408__B _05112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15953_ net1403 vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__inv_2
XANTENNA__09605__C net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10027_ net561 net552 net534 vssd1 vssd1 vccd1 vccd1 _06367_ sky130_fd_sc_hd__or3_1
X_14904_ net1213 vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_129_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15884_ net1360 vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__inv_2
XANTENNA__10142__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17623_ clknet_leaf_5_wb_clk_i _03308_ _01564_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14835_ net1419 vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_125_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11643__S net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17554_ clknet_leaf_144_wb_clk_i _03241_ _01537_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11978_ net2739 net256 net471 vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__mux2_1
X_14766_ net1293 vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__inv_2
XANTENNA__13092__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09835__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08518__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16505_ clknet_leaf_2_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[3\]
+ _00488_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13717_ team_01_WB.instance_to_wrap.cpu.c0.count\[7\] _04103_ net2890 vssd1 vssd1
+ vccd1 vccd1 _04128_ sky130_fd_sc_hd__a21oi_1
X_10929_ net563 _07253_ _07264_ _07268_ vssd1 vssd1 vccd1 vccd1 _07269_ sky130_fd_sc_hd__a211o_2
X_14697_ net1195 vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__inv_2
X_17485_ clknet_leaf_108_wb_clk_i _03172_ _01468_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16436_ clknet_leaf_133_wb_clk_i _02190_ _00419_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13648_ net187 _04081_ _04082_ net728 vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__a211o_1
XFILLER_0_73_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12474__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16367_ clknet_leaf_91_wb_clk_i net2953 _00350_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[90\]
+ sky130_fd_sc_hd__dfrtp_1
X_13579_ _03917_ _04024_ vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__nor2_1
XANTENNA__14255__A net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15318_ net1247 vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__inv_2
XANTENNA__08271__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16298_ clknet_leaf_100_wb_clk_i _02052_ _00281_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[21\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_112_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13147__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15249_ net1420 vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__inv_2
XANTENNA__11158__A1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09810_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[14\] net816 net746 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06150_ sky130_fd_sc_hd__a22o_1
Xfanout307 _07935_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__buf_2
XANTENNA__11818__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10905__B2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11169__C_N _07308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout318 net320 vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__buf_2
XANTENNA__10381__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13304__C1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09741_ net1132 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[20\] net957
+ vssd1 vssd1 vccd1 vccd1 _06081_ sky130_fd_sc_hd__and3_1
XANTENNA__15814__A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09672_ net1136 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[22\] net956
+ vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__and3_1
XANTENNA__10764__S0 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08623_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[11\] net683 _04962_
+ net705 vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__a211o_1
XANTENNA__12649__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08554_ net1077 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[19\] net906
+ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_85_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16418__Q team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08485_ net1100 net941 vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__and2_2
XANTENNA__08495__D1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11633__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout434_A _07964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10841__A0 _06065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14032__B1 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12892__B net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout601_A _04754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12384__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1343_A net1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09106_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[13\] net667 _05427_ _05438_
+ _05441_ vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_131_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09037_ _05006_ _05338_ _05374_ vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__and3_1
XANTENNA__11301__B _05153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1131_X net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1229_X net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold350 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1885 sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1896 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08450__X _04790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12897__A1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout970_A _04645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout689_X net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold372 _01927_ vssd1 vssd1 vccd1 vccd1 net1907 sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1918 sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1929 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14099__B1 _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout830 net831 vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__clkbuf_2
Xfanout841 net842 vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__clkbuf_2
Xfanout852 net853 vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__clkbuf_4
X_09939_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[4\] net764 net623 vssd1
+ vssd1 vccd1 vccd1 _06279_ sky130_fd_sc_hd__o21a_1
Xfanout863 net864 vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__clkbuf_4
Xfanout874 net876 vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__clkbuf_2
Xfanout885 net886 vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__buf_2
Xfanout896 net897 vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__buf_4
X_12950_ net1038 net585 _03709_ vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__a21oi_2
XANTENNA__11321__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10124__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1050 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[38\] vssd1 vssd1 vccd1 vccd1
+ net2585 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1061 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2596 sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ net2285 net205 net479 vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__mux2_1
Xhold1072 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2607 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1083 team_01_WB.instance_to_wrap.cpu.f0.num\[22\] vssd1 vssd1 vccd1 vccd1 net2618
+ sky130_fd_sc_hd__dlygate4sd3_1
X_12881_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[28\] _03661_ net1036 vssd1
+ vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1094 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[54\] vssd1 vssd1 vccd1 vccd1
+ net2629 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12559__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14620_ net1309 vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__inv_2
X_11832_ net2009 net246 net489 vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__mux2_1
XANTENNA__10220__X _06560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09278__B1 _05617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14551_ net1406 vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__inv_2
XANTENNA__09160__C net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11763_ net2261 net210 net495 vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_155_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12821__B2 _03643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ net554 _06928_ vssd1 vssd1 vccd1 vccd1 _07054_ sky130_fd_sc_hd__and2_2
X_13502_ net720 _07019_ net1073 vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_120_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ net1356 vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__inv_2
X_17270_ clknet_leaf_24_wb_clk_i _02957_ _01253_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11694_ net1890 net253 net499 vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__mux2_1
XANTENNA__14023__B1 _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16221_ clknet_leaf_130_wb_clk_i net1648 _00209_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__dfrtp_1
X_13433_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\] net595 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\]
+ vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__a21oi_1
X_10645_ net507 net505 net543 vssd1 vssd1 vccd1 vccd1 _06985_ sky130_fd_sc_hd__mux2_1
XANTENNA__12294__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16152_ clknet_leaf_131_wb_clk_i _01915_ _00140_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13364_ net1070 net1071 vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10576_ net503 _06882_ net369 vssd1 vssd1 vccd1 vccd1 _06916_ sky130_fd_sc_hd__o21a_1
XFILLER_0_63_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09450__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12315_ net2458 net301 net432 vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15103_ net1317 vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__inv_2
X_16083_ clknet_leaf_131_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[5\]
+ _00071_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13295_ _03751_ _03780_ _04621_ vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10890__X _07230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13534__C1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15034_ net1372 vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__inv_2
X_12246_ net2343 net225 net439 vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08801__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_91_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_82_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12177_ net3147 net284 net449 vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__mux2_1
XANTENNA__10542__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_20_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10363__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11128_ net525 _07256_ _07467_ _06906_ vssd1 vssd1 vccd1 vccd1 _07468_ sky130_fd_sc_hd__o22ai_1
X_16985_ clknet_leaf_103_wb_clk_i _02672_ _00968_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11059_ net555 _06281_ _07384_ _06251_ _05076_ vssd1 vssd1 vccd1 vccd1 _07399_ sky130_fd_sc_hd__a32o_1
X_15936_ net1402 vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__inv_2
XANTENNA__18010__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10115__A2 _04636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09632__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15867_ net1202 vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__inv_2
XANTENNA__12469__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11226__X _07566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17606_ clknet_leaf_86_wb_clk_i _03293_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_14818_ net1320 vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09269__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15798_ net1232 vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_103_Left_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16238__Q net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17537_ clknet_leaf_53_wb_clk_i _03224_ _01520_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_14749_ net1187 vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__inv_2
XANTENNA__12812__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08270_ net2847 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[3\] net1055 vssd1 vssd1
+ vccd1 vccd1 _03417_ sky130_fd_sc_hd__mux2_1
X_17468_ clknet_leaf_60_wb_clk_i _03155_ _01451_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_2__f_wb_clk_i_X clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16419_ clknet_leaf_138_wb_clk_i _02173_ _00402_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13368__A2 _04579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17399_ clknet_leaf_14_wb_clk_i _03086_ _01382_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09441__A0 _05779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10354__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07985_ team_01_WB.instance_to_wrap.cpu.f0.i\[10\] vssd1 vssd1 vccd1 vccd1 _04483_
+ sky130_fd_sc_hd__inv_2
XANTENNA_fanout384_A _03570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09724_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[21\] net765 net624 vssd1
+ vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_87_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10106__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09542__A net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09655_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[23\] net763 net622 vssd1
+ vssd1 vccd1 vccd1 _05995_ sky130_fd_sc_hd__o21a_1
XANTENNA__12379__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1293_A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout649_A _04823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08606_ net1168 _04846_ _04845_ vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__a21o_1
XANTENNA__11136__X _07476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09586_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[25\] net785 net761 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__a22o_1
X_08537_ _04873_ _04874_ _04875_ _04876_ vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__nor4_1
XANTENNA_fanout816_A _04636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout437_X net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10814__B1 _07153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08468_ net1024 net902 vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__and2_2
XFILLER_0_92_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14005__B1 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08445__X _04785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout604_X net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08399_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\] net710 net621 _04724_ vssd1
+ vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__a22oi_2
XTAP_TAPCELL_ROW_150_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10430_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[27\] net811 _06757_ _06760_
+ _06761_ vssd1 vssd1 vccd1 vccd1 _06770_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_104_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09432__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08324__C net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10361_ _06683_ _06698_ _06699_ _06700_ vssd1 vssd1 vccd1 vccd1 _06701_ sky130_fd_sc_hd__or4_1
XFILLER_0_115_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12842__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12100_ net3124 net203 net455 vssd1 vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13516__C1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13080_ net2987 net2620 net853 vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10292_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[19\] net734 _06629_ _06630_
+ _06631_ vssd1 vssd1 vccd1 vccd1 _06632_ sky130_fd_sc_hd__a2111o_1
XANTENNA__17707__Q team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout973_X net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12031_ net2581 net245 net465 vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__mux2_1
XANTENNA__08538__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold180 net98 vssd1 vssd1 vccd1 vccd1 net1715 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold191 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[11\] vssd1 vssd1 vccd1 vccd1
+ net1726 sky130_fd_sc_hd__dlygate4sd3_1
X_17954__1469 vssd1 vssd1 vccd1 vccd1 _17954__1469/HI net1469 sky130_fd_sc_hd__conb_1
XANTENNA__08340__B net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout660 net661 vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11166__A2_N _07499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout671 _04797_ vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__buf_8
X_16770_ clknet_leaf_76_wb_clk_i _02457_ _00753_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout682 net683 vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__clkbuf_8
Xfanout693 _04771_ vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__buf_8
X_13982_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[104\] _04252_ _04268_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[72\]
+ vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__a22o_1
XANTENNA__08994__C net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15721_ net1296 vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__inv_2
X_12933_ net356 _03697_ _03698_ net869 net3158 vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__a32o_1
XANTENNA__12289__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15652_ net1220 vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_122_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13405__C net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12864_ net2978 net313 net380 vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__mux2_1
XANTENNA__16058__Q team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14603_ net1357 vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__inv_2
X_11815_ net2807 net301 net492 vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12795_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[11\] _07207_ net1035 vssd1 vssd1
+ vccd1 vccd1 _03625_ sky130_fd_sc_hd__mux2_1
X_15583_ net1315 vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11921__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17322_ clknet_leaf_33_wb_clk_i _03009_ _01305_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11746_ _07932_ _07933_ _07934_ net613 vssd1 vssd1 vccd1 vccd1 _07935_ sky130_fd_sc_hd__a22o_4
X_14534_ net1351 vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17253_ clknet_leaf_51_wb_clk_i _02940_ _01236_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11677_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] _07811_ vssd1 vssd1
+ vccd1 vccd1 _07879_ sky130_fd_sc_hd__xnor2_1
X_14465_ net1188 vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16204_ clknet_leaf_133_wb_clk_i _01964_ _00192_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10628_ _04706_ net503 net543 vssd1 vssd1 vccd1 vccd1 _06968_ sky130_fd_sc_hd__mux2_1
X_13416_ _03871_ _03876_ _03870_ vssd1 vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__a21o_1
X_17184_ clknet_leaf_46_wb_clk_i _02871_ _01167_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_14396_ net1188 vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__inv_2
XANTENNA__09423__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11230__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16135_ clknet_leaf_157_wb_clk_i _00009_ _00123_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.curr_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13347_ net586 _07687_ _03820_ net829 vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__a31o_1
X_10559_ net542 _06896_ _06898_ vssd1 vssd1 vccd1 vccd1 _06899_ sky130_fd_sc_hd__o21a_1
XFILLER_0_12_728 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_106_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16066_ clknet_leaf_155_wb_clk_i _01859_ _00054_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\]
+ sky130_fd_sc_hd__dfrtp_4
X_13278_ _03748_ _03766_ _04518_ vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__a21oi_1
X_15017_ net1295 vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__inv_2
XANTENNA__13522__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12229_ net2557 net214 net441 vssd1 vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__mux2_1
XANTENNA__11595__C team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11533__B2 net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16968_ clknet_leaf_63_wb_clk_i _02655_ _00951_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13286__B2 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10004__C net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15919_ net1412 vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__inv_2
XANTENNA__12199__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16899_ clknet_leaf_23_wb_clk_i _02586_ _00882_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_09440_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\] net710 net594 vssd1 vssd1
+ vccd1 vccd1 _05780_ sky130_fd_sc_hd__a21o_1
XANTENNA__08701__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12921__B1_N net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13589__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08409__C _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09371_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[26\] net694 net691 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10795__X _07135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11831__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08322_ net1161 net1165 net1166 net1158 vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__and4b_4
XANTENNA_clkbuf_leaf_58_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_24_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08706__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10955__B _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08253_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[28\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[20\]
+ net1045 vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11132__A net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13746__C1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08184_ net2457 net2815 net1056 vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09414__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08768__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12662__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1041_A team_01_WB.instance_to_wrap.cpu.RU0.InstrRead vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1139_A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11772__A1 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09537__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13513__A2 _07088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10327__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11524__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1306_A net1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout766_A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout387_X net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07968_ team_01_WB.instance_to_wrap.cpu.f0.i\[29\] vssd1 vssd1 vccd1 vccd1 _04466_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_96_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09707_ net1154 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[21\] net949
+ vssd1 vssd1 vccd1 vccd1 _06047_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_143_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout554_X net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_97_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09703__C net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09638_ net993 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[23\] net956 vssd1
+ vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__and3_1
XANTENNA__11026__B net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout721_X net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09569_ net1149 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[25\] net979
+ vssd1 vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__and3_1
XANTENNA__12837__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout819_X net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11600_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\]
+ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] _07814_ vssd1 vssd1 vccd1 vccd1
+ _07817_ sky130_fd_sc_hd__and4_1
XANTENNA__12788__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12580_ net2014 net278 net399 vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11531_ net2518 net1171 net588 net1121 vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__a22o_1
XANTENNA__11460__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08335__B net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14250_ net1226 vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__inv_2
XANTENNA__14056__C _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11462_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[7\] _07757_ net877 vssd1 vssd1
+ vccd1 vccd1 _07758_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_52_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09405__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13201_ net7 net837 _03738_ net2178 vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10413_ net1132 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[27\] net972
+ vssd1 vssd1 vccd1 vccd1 _06753_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_78_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14181_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[11\] _04452_ vssd1 vssd1 vccd1
+ vccd1 _04453_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_78_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11393_ _04466_ _07715_ _07719_ net323 vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__o211a_1
XANTENNA__12572__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13132_ net77 net844 net632 net1634 vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__a22o_1
XANTENNA__08989__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10344_ net1139 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[17\] net984
+ vssd1 vssd1 vccd1 vccd1 _06684_ sky130_fd_sc_hd__and3_1
XANTENNA_input62_A wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13063_ net2854 net2769 net857 vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__mux2_1
X_17940_ net1455 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
X_10275_ net990 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[19\] net954 vssd1
+ vssd1 vccd1 vccd1 _06615_ sky130_fd_sc_hd__and3_1
XANTENNA__11515__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12014_ net2531 net249 net469 vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__mux2_1
Xfanout1400 net1409 vssd1 vssd1 vccd1 vccd1 net1400 sky130_fd_sc_hd__buf_4
Xfanout1411 net1414 vssd1 vssd1 vccd1 vccd1 net1411 sky130_fd_sc_hd__buf_4
Xfanout1422 net1425 vssd1 vssd1 vccd1 vccd1 net1422 sky130_fd_sc_hd__buf_2
X_17871_ clknet_leaf_138_wb_clk_i _03546_ _01811_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11916__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16822_ clknet_leaf_29_wb_clk_i _02509_ _00805_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout490 _07947_ vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__buf_4
X_16753_ clknet_leaf_113_wb_clk_i _02440_ _00736_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13965_ _04219_ _04231_ vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__nand2_2
X_15704_ net1223 vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12916_ net356 _03685_ _03686_ net869 net1557 vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__a32o_1
X_16684_ clknet_leaf_16_wb_clk_i _02371_ _00667_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13896_ _04141_ net572 _04199_ vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__and3b_1
XFILLER_0_76_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15635_ net1419 vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12747__S net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14087__X _04375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12847_ net2019 net235 net379 vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11651__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12779__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13432__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15566_ net1300 vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12778_ net362 _03612_ _03613_ net1061 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\]
+ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__a32o_1
XANTENNA__09644__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17305_ clknet_leaf_104_wb_clk_i _02992_ _01288_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14517_ net1412 vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__inv_2
X_11729_ net613 _07799_ _07920_ _07919_ vssd1 vssd1 vccd1 vccd1 _07921_ sky130_fd_sc_hd__a31o_4
X_15497_ net1294 vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10494__C net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17236_ clknet_leaf_66_wb_clk_i _02923_ _01219_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14448_ net1305 vssd1 vssd1 vccd1 vccd1 _00242_ sky130_fd_sc_hd__inv_2
XANTENNA__08813__X _05153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12482__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17167_ clknet_leaf_31_wb_clk_i _02854_ _01150_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold905 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[34\] vssd1 vssd1 vccd1 vccd1
+ net2440 sky130_fd_sc_hd__dlygate4sd3_1
X_14379_ net1195 vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__inv_2
Xhold916 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2451 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11754__A1 _07438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold927 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2462 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08899__C net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16118_ clknet_leaf_136_wb_clk_i _01893_ _00106_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[25\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold938 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17098_ clknet_leaf_32_wb_clk_i _02785_ _01081_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold949 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2484 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08940_ net1112 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[6\] net927 vssd1
+ vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__and3_1
X_16049_ clknet_leaf_148_wb_clk_i _01842_ _00037_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_08871_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[3\] _04800_ net651 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[3\]
+ _05196_ vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_131_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1605 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3140 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1616 team_01_WB.instance_to_wrap.cpu.c0.count\[11\] vssd1 vssd1 vccd1 vccd1 net3151
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1627 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net3162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1638 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 net3173
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1649 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 net3184
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_35_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09423_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[28\] net682 net678 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__a22o_1
XANTENNA__12657__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09354_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[25\] net699 net649 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1089_A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08436__A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17953__1468 vssd1 vssd1 vccd1 vccd1 _17953__1468/HI net1468 sky130_fd_sc_hd__conb_1
XFILLER_0_19_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08305_ net1159 net1164 net1168 net1162 vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09285_ net1084 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[22\] net887
+ vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__and3_1
XANTENNA__13982__A2 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout514_A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1256_A net1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08236_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[45\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[37\]
+ net1051 vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13195__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08167_ net2350 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[106\] net1052 vssd1 vssd1
+ vccd1 vccd1 _03520_ sky130_fd_sc_hd__mux2_1
XANTENNA__13734__A2 _04516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12392__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12942__B1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08098_ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[4\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[7\]
+ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[6\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__or4b_1
XANTENNA_fanout883_A _04803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1531_A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[22\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10206__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_148_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_148_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_145_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10060_ _06367_ _06368_ _06366_ vssd1 vssd1 vccd1 vccd1 _06400_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_145_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout671_X net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout769_X net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11736__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout936_X net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15732__A net1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13750_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[0\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__nand2_1
X_10962_ net539 _07301_ vssd1 vssd1 vccd1 vccd1 _07302_ sky130_fd_sc_hd__nand2_1
XANTENNA__09874__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09730__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12701_ net1917 net236 net383 vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__mux2_1
XANTENNA__11681__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10893_ _06677_ _07113_ net343 vssd1 vssd1 vccd1 vccd1 _07233_ sky130_fd_sc_hd__a21oi_1
X_13681_ team_01_WB.instance_to_wrap.cpu.c0.count\[7\] _04103_ vssd1 vssd1 vccd1 vccd1
+ _04104_ sky130_fd_sc_hd__nand2_1
XANTENNA__12567__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15420_ net1246 vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__inv_2
X_12632_ net1937 net242 net392 vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__mux2_1
XANTENNA__08346__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10595__B _06902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12563_ net3130 net272 net401 vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__mux2_1
X_15351_ net1244 vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14302_ net1328 vssd1 vssd1 vccd1 vccd1 _00096_ sky130_fd_sc_hd__inv_2
XANTENNA__09876__S net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11514_ net1555 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[4\] net877 vssd1 vssd1
+ vccd1 vccd1 _03335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15282_ net1266 vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_117_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12494_ net3022 net210 net407 vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_117_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17021_ clknet_leaf_58_wb_clk_i _02708_ _01004_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13186__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15179__A net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14233_ net1308 vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__inv_2
X_11445_ team_01_WB.instance_to_wrap.cpu.f0.i\[4\] _07674_ net325 vssd1 vssd1 vccd1
+ vccd1 _07747_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11197__C1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10539__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12933__B1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14164_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[4\] _04188_ vssd1 vssd1 vccd1
+ vccd1 _04443_ sky130_fd_sc_hd__xnor2_1
X_11376_ _04477_ _07704_ vssd1 vssd1 vccd1 vccd1 _07705_ sky130_fd_sc_hd__nor2_1
XANTENNA__09608__C net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16071__Q team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08512__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_156_Right_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13115_ net1573 net844 net633 team_01_WB.instance_to_wrap.a1.ADR_I\[28\] vssd1 vssd1
+ vccd1 vccd1 _02026_ sky130_fd_sc_hd__a22o_1
X_10327_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[18\] net794 _06664_ _06665_
+ _06666_ vssd1 vssd1 vccd1 vccd1 _06667_ sky130_fd_sc_hd__a2111o_1
X_14095_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[29\] _04243_ _04252_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[109\]
+ _04381_ vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__a221o_1
X_17923_ net1530 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
X_13046_ net2388 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[48\] net857 vssd1 vssd1
+ vccd1 vccd1 _02079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10258_ _06221_ _06469_ _06472_ _06597_ vssd1 vssd1 vccd1 vccd1 _06598_ sky130_fd_sc_hd__or4_2
XANTENNA__11646__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08365__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1230 net1232 vssd1 vssd1 vccd1 vccd1 net1230 sky130_fd_sc_hd__buf_4
XANTENNA__13427__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1241 net1242 vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__buf_2
X_17854_ clknet_leaf_98_wb_clk_i _03530_ _01794_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[124\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__10172__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10189_ _04750_ _05376_ _05006_ vssd1 vssd1 vccd1 vccd1 _06529_ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1252 net1303 vssd1 vssd1 vccd1 vccd1 net1252 sky130_fd_sc_hd__buf_2
Xfanout1263 net1264 vssd1 vssd1 vccd1 vccd1 net1263 sky130_fd_sc_hd__buf_2
Xfanout1274 net1275 vssd1 vssd1 vccd1 vccd1 net1274 sky130_fd_sc_hd__buf_4
X_16805_ clknet_leaf_51_wb_clk_i _02492_ _00788_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1285 net1302 vssd1 vssd1 vccd1 vccd1 net1285 sky130_fd_sc_hd__buf_2
Xfanout1296 net1301 vssd1 vssd1 vccd1 vccd1 net1296 sky130_fd_sc_hd__buf_2
XANTENNA__09343__C net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17785_ clknet_leaf_121_wb_clk_i _03461_ _01725_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[55\]
+ sky130_fd_sc_hd__dfrtp_1
X_14997_ net1276 vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16736_ clknet_leaf_48_wb_clk_i _02423_ _00719_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13948_ _04227_ _04237_ _04239_ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__and3_4
XANTENNA__09865__B1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09640__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12477__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16667_ clknet_leaf_68_wb_clk_i _02354_ _00650_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17630__Q team_01_WB.instance_to_wrap.cpu.IG0.Instr\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13879_ team_01_WB.instance_to_wrap.cpu.RU0.state\[0\] _03575_ _04136_ _00005_ vssd1
+ vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_read_i sky130_fd_sc_hd__a31o_1
XFILLER_0_8_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15618_ net1351 vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16598_ clknet_leaf_15_wb_clk_i _02285_ _00581_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[30\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_72_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15549_ net1313 vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__inv_2
X_09070_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[12\] net661 _05387_
+ _05399_ _05402_ vssd1 vssd1 vccd1 vccd1 _05410_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_21_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08021_ _04505_ _04516_ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__nor2_1
X_17219_ clknet_leaf_66_wb_clk_i _02906_ _01202_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10725__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11727__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11410__A team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12924__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold702 _03505_ vssd1 vssd1 vccd1 vccd1 net2237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold724 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2259 sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2270 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold746 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[9\] vssd1 vssd1 vccd1 vccd1 net2281
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold757 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2303 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold779 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2314 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09972_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[3\] net765 net624 vssd1
+ vssd1 vccd1 vccd1 _06312_ sky130_fd_sc_hd__o21a_1
XANTENNA__09148__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08923_ net525 net516 vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__nand2_4
XANTENNA__14141__A2 _04230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08356__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout297_A _07921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1402 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2937 sky130_fd_sc_hd__dlygate4sd3_1
X_08854_ net1106 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[3\] net907 vssd1
+ vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__and3_1
Xhold1413 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2948 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10163__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1424 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2959 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1004_A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1435 team_01_WB.instance_to_wrap.cpu.f0.num\[20\] vssd1 vssd1 vccd1 vccd1 net2970
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1446 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2981 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08785_ net1014 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[0\] net910 vssd1
+ vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__and3_1
Xhold1457 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[98\] vssd1 vssd1 vccd1 vccd1
+ net2992 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_140_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1468 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net3003 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout464_A _07954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1479 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[10\] vssd1 vssd1 vccd1 vccd1 net3014
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09856__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13652__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12387__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11663__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout631_A _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1373_A net1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09406_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[27\] net687 net671 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[27\]
+ _05745_ vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_66_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09337_ _05661_ _05674_ _05675_ _05676_ vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_138_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10983__X _07323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09268_ net1080 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[20\] net906
+ net656 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[20\] vssd1 vssd1 vccd1
+ vccd1 _05608_ sky130_fd_sc_hd__a32o_1
XANTENNA__08453__X _04793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08219_ net2725 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[54\] net1043 vssd1 vssd1
+ vccd1 vccd1 _03468_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09199_ net1082 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[17\] net900
+ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1426_X net1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11230_ _05934_ _05965_ _07568_ net343 vssd1 vssd1 vccd1 vccd1 _07570_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_112_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11161_ _05076_ net332 _07500_ net370 vssd1 vssd1 vccd1 vccd1 _07501_ sky130_fd_sc_hd__a211oi_1
XANTENNA__12850__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10112_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[6\] net753 net750 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06452_ sky130_fd_sc_hd__a22o_1
XANTENNA__14132__A2 _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11092_ net534 _06366_ vssd1 vssd1 vccd1 vccd1 _07432_ sky130_fd_sc_hd__nor2_1
X_10043_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[0\] net817 net791 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06383_ sky130_fd_sc_hd__a22o_1
X_14920_ net1375 vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__inv_2
Xhold40 net79 vssd1 vssd1 vccd1 vccd1 net1575 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 _02022_ vssd1 vssd1 vccd1 vccd1 net1586 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 _02025_ vssd1 vssd1 vccd1 vccd1 net1597 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input25_A DAT_I[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold73 _02010_ vssd1 vssd1 vccd1 vccd1 net1608 sky130_fd_sc_hd__dlygate4sd3_1
X_14851_ net1221 vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__inv_2
Xhold84 _01988_ vssd1 vssd1 vccd1 vccd1 net1619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 team_01_WB.instance_to_wrap.a1.ADR_I\[10\] vssd1 vssd1 vccd1 vccd1 net1630
+ sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ _01836_ _04164_ _04173_ _01837_ vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__a31o_1
X_17570_ clknet_leaf_86_wb_clk_i _03257_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13643__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14782_ net1316 vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__inv_2
X_11994_ net2045 net222 net467 vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__mux2_1
XANTENNA__08628__X _04968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09311__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16521_ clknet_leaf_0_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[19\]
+ _00504_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13733_ team_01_WB.instance_to_wrap.cpu.DM0.dhit team_01_WB.instance_to_wrap.cpu.f0.state\[3\]
+ team_01_WB.instance_to_wrap.cpu.f0.state\[0\] team_01_WB.EN_VAL_REG vssd1 vssd1
+ vccd1 vccd1 _04134_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10945_ _06129_ _06158_ _06188_ _06216_ net550 net539 vssd1 vssd1 vccd1 vccd1 _07285_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12297__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_45_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_128_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16452_ clknet_leaf_106_wb_clk_i _02206_ _00435_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13664_ net722 _07489_ net1075 vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__o21a_1
X_10876_ net524 _07215_ _07213_ vssd1 vssd1 vccd1 vccd1 _07216_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_39_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15403_ net1397 vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__inv_2
XANTENNA__16066__Q team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12615_ net2409 net293 net397 vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__mux2_1
XANTENNA__11214__B _07207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16383_ clknet_leaf_90_wb_clk_i net2773 _00366_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13595_ net187 _04037_ _04038_ net726 vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__a211o_1
XFILLER_0_155_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15334_ net1405 vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__inv_2
X_12546_ net1930 net300 net406 vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13159__B1 _03734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15265_ net1278 vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12477_ net2528 net228 net411 vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_4 _03654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12906__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17004_ clknet_leaf_19_wb_clk_i _02691_ _00987_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_14216_ net1910 vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11428_ _07679_ _07700_ team_01_WB.instance_to_wrap.cpu.f0.i\[13\] vssd1 vssd1 vccd1
+ vccd1 _07739_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15196_ net1244 vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11359_ net1071 _07681_ vssd1 vssd1 vccd1 vccd1 _07688_ sky130_fd_sc_hd__nand2_1
X_14147_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[39\] _04221_ _04233_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[71\]
+ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__a22o_1
XANTENNA__10393__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09635__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14123__A2 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14078_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[52\] _04236_ _04250_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[124\]
+ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__a22o_1
X_17952__1467 vssd1 vssd1 vccd1 vccd1 _17952__1467/HI net1467 sky130_fd_sc_hd__conb_1
X_17906_ net1441 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
X_13029_ net2597 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[65\] net865 vssd1 vssd1
+ vccd1 vccd1 _02096_ sky130_fd_sc_hd__mux2_1
Xfanout1060 net1061 vssd1 vssd1 vccd1 vccd1 net1060 sky130_fd_sc_hd__clkbuf_4
Xfanout1071 net1072 vssd1 vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__buf_2
X_17837_ clknet_leaf_95_wb_clk_i _03513_ _01777_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[107\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09550__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1082 net1089 vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__clkbuf_2
Xfanout1093 net1096 vssd1 vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_156_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08570_ net999 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[19\] net883 vssd1
+ vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17768_ clknet_leaf_117_wb_clk_i _03444_ _01708_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13634__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16719_ clknet_leaf_31_wb_clk_i _02406_ _00702_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17699_ clknet_leaf_134_wb_clk_i _03383_ _01640_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_18_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12000__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09122_ net1022 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[14\] net889 vssd1
+ vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08714__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09053_ net1029 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[12\] net912
+ vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_40_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout212_A net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08433__B _04770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08004_ net1682 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[0\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_142_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09369__A2 _04766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold510 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2045 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold521 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2056 sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2067 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13570__B1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold543 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2078 sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2089 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12670__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold565 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2100 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08041__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10384__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold576 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2111 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1219_A net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold587 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2133 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14114__A2 _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09955_ net1155 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[3\] net980 vssd1
+ vssd1 vccd1 vccd1 _06295_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout679_A _04789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08906_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[2\] net931 vssd1
+ vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__and3_1
XANTENNA__10136__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09886_ net998 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[5\] net964 vssd1
+ vssd1 vccd1 vccd1 _06226_ sky130_fd_sc_hd__and3_1
Xhold1210 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[97\] vssd1 vssd1 vccd1 vccd1
+ net2745 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1221 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[79\] vssd1 vssd1 vccd1 vccd1
+ net2756 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1232 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[56\] vssd1 vssd1 vccd1 vccd1
+ net2767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1243 team_01_WB.instance_to_wrap.cpu.K0.count\[1\] vssd1 vssd1 vccd1 vccd1 net2778
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08837_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[1\] net669 net668 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__a22o_1
Xhold1254 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 net2789
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout846_A net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout467_X net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1265 _03495_ vssd1 vssd1 vccd1 vccd1 net2800 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1276 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2811 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1287 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2822 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09829__B1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08768_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[4\] net697 _05079_ _05083_
+ _05097_ vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08448__X _04788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1298 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2833 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08699_ _05030_ _05031_ _05037_ _05038_ vssd1 vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__or4_2
XFILLER_0_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08501__B1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13006__S net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10730_ net553 _07069_ vssd1 vssd1 vccd1 vccd1 _07070_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_64_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11034__B net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10661_ _06438_ _06562_ net552 vssd1 vssd1 vccd1 vccd1 _07001_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout801_X net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12845__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11939__A1 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12400_ net1925 net202 net420 vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_149_Left_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13380_ _03839_ _03840_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10592_ net523 _06894_ _06906_ _06909_ vssd1 vssd1 vccd1 vccd1 _06932_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_134_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_153_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12331_ net3079 net206 net429 vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15050_ net1385 vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__inv_2
X_12262_ net2473 net215 net435 vssd1 vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09158__C net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14001_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[9\] _04226_ _04254_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[97\]
+ vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__a22o_1
X_11213_ net562 _07543_ _07544_ _07552_ vssd1 vssd1 vccd1 vccd1 _07553_ sky130_fd_sc_hd__a31o_2
XFILLER_0_142_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12580__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12193_ net2463 net218 net445 vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__mux2_1
XANTENNA__08630__Y _04970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10914__A2 _06526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11144_ _07327_ _07329_ net535 vssd1 vssd1 vccd1 vccd1 _07484_ sky130_fd_sc_hd__mux2_1
XANTENNA__14105__A2 _04221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09780__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__buf_2
XFILLER_0_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__buf_2
X_11075_ _07413_ _07414_ _07359_ vssd1 vssd1 vccd1 vccd1 _07415_ sky130_fd_sc_hd__a21oi_1
X_15952_ net1402 vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__inv_2
X_10026_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] _06365_ _04628_ vssd1
+ vssd1 vccd1 vccd1 _06366_ sky130_fd_sc_hd__mux2_2
X_14903_ net1243 vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_129_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15883_ net1347 vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_129_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11924__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17622_ clknet_leaf_5_wb_clk_i _03307_ _01563_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_14834_ net1291 vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__inv_2
XANTENNA__13616__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11627__A0 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17553_ clknet_leaf_113_wb_clk_i _03240_ _01536_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_14765_ net1262 vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__inv_2
X_11977_ net2817 net259 net473 vssd1 vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16504_ clknet_leaf_2_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[2\]
+ _00487_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13716_ _04103_ _04127_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[6\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_156_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10928_ net553 _07267_ vssd1 vssd1 vccd1 vccd1 _07268_ sky130_fd_sc_hd__nor2_1
X_17484_ clknet_leaf_149_wb_clk_i _03171_ _01467_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_14696_ net1198 vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16435_ clknet_leaf_132_wb_clk_i _02189_ _00418_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13647_ net198 net194 _07925_ net644 vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10859_ _06129_ _06707_ net371 _06671_ net533 net544 vssd1 vssd1 vccd1 vccd1 _07199_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_2_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13440__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16366_ clknet_leaf_87_wb_clk_i _02120_ _00349_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[89\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13578_ _03914_ _03916_ vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__nor2_1
X_15317_ net1287 vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12529_ net2982 net207 net404 vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16297_ clknet_leaf_118_wb_clk_i _02051_ _00280_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[20\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_83_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15248_ net1271 vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12490__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15179_ net1397 vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__inv_2
XANTENNA__10905__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout308 _07935_ vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__buf_1
XFILLER_0_10_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09771__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout319 net320 vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__clkbuf_2
X_09740_ net1145 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[20\] net959
+ vssd1 vssd1 vccd1 vccd1 _06080_ sky130_fd_sc_hd__and3_1
XANTENNA__10118__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
.ends

